magic
tech scmos
timestamp 1758851824
<< nwell >>
rect -47 0 41 20
<< pwell >>
rect -47 -30 41 0
rect -47 -31 40 -30
<< ntransistor >>
rect -32 -11 -27 -6
rect -7 -11 -3 -6
rect 1 -11 5 -6
rect 12 -11 16 -6
rect 20 -11 24 -6
<< ptransistor >>
rect -32 6 -27 11
rect -7 6 -3 11
rect 1 6 5 11
rect 12 6 16 11
rect 20 6 24 11
<< ndiffusion >>
rect -36 -11 -32 -6
rect -27 -11 -24 -6
rect -15 -11 -14 -6
rect -9 -11 -7 -6
rect -3 -11 1 -6
rect 5 -11 6 -6
rect 11 -11 12 -6
rect 16 -11 20 -6
rect 24 -11 29 -6
rect 34 -11 35 -6
<< pdiffusion >>
rect -36 6 -32 11
rect -27 6 -24 11
rect -15 6 -14 11
rect -9 6 -7 11
rect -3 6 1 11
rect 5 6 6 11
rect 11 6 12 11
rect 16 6 20 11
rect 24 6 29 11
rect 34 6 35 11
<< ndcontact >>
rect -41 -11 -36 -6
rect -24 -11 -19 -6
rect -14 -11 -9 -6
rect 6 -11 11 -6
rect 29 -11 34 -6
<< pdcontact >>
rect -41 6 -36 11
rect -24 6 -19 11
rect -14 6 -9 11
rect 6 6 11 11
rect 29 6 34 11
<< polysilicon >>
rect -32 11 -27 15
rect -7 11 -3 16
rect 1 11 5 14
rect 12 11 16 14
rect 20 11 24 16
rect -32 3 -27 6
rect -32 -6 -27 -2
rect -7 -6 -3 6
rect 1 2 5 6
rect 12 2 16 6
rect 1 -6 5 -2
rect 12 -6 16 -2
rect 20 -6 24 6
rect -32 -17 -27 -11
rect -7 -24 -3 -11
rect 1 -14 5 -11
rect 12 -17 16 -11
rect 20 -18 24 -11
<< polycontact >>
rect 1 14 6 19
rect 11 14 16 19
rect -32 -2 -27 3
rect 1 -19 6 -14
rect 11 -22 16 -17
rect 20 -23 25 -18
rect -8 -29 -3 -24
<< metal1 >>
rect 11 19 41 20
rect -30 16 1 19
rect -42 11 -35 12
rect -42 6 -41 11
rect -36 6 -35 11
rect -42 5 -35 6
rect -30 3 -27 16
rect 16 17 41 19
rect -15 11 -8 12
rect 28 11 35 12
rect -42 -6 -35 -5
rect -42 -11 -41 -6
rect -36 -11 -35 -6
rect -42 -12 -35 -11
rect -30 -16 -27 -2
rect -22 -6 -19 6
rect -15 6 -14 11
rect -9 6 -8 11
rect -15 5 -8 6
rect 7 0 11 6
rect 28 6 29 11
rect 34 6 35 11
rect 28 5 35 6
rect 16 0 23 3
rect 7 -3 23 0
rect -22 -15 -19 -11
rect -15 -6 -8 -5
rect 7 -6 11 -3
rect 16 -4 23 -3
rect -15 -11 -14 -6
rect -9 -11 -8 -6
rect 28 -6 35 -5
rect 28 -11 29 -6
rect 34 -11 35 -6
rect -15 -12 -8 -11
rect 28 -12 35 -11
rect -33 -23 -26 -16
rect -22 -18 1 -15
rect -9 -29 -8 -24
rect 3 -27 6 -19
rect 10 -17 17 -16
rect 10 -22 11 -17
rect 16 -22 17 -17
rect 10 -23 17 -22
rect 38 -27 41 17
rect 3 -30 41 -27
<< metal2 >>
rect -42 11 -35 12
rect -15 11 -8 12
rect 28 11 35 12
rect -42 7 35 11
rect -42 6 11 7
rect -42 5 -35 6
rect -15 5 -8 6
rect 28 5 35 7
rect 16 -4 23 3
rect -42 -6 -35 -5
rect -15 -6 -8 -5
rect -42 -8 11 -6
rect 28 -8 35 -5
rect -42 -11 35 -8
rect -42 -12 -35 -11
rect -15 -12 -8 -11
rect 28 -12 35 -11
rect -33 -17 -26 -16
rect 10 -17 17 -16
rect -33 -21 17 -17
rect -33 -23 -26 -21
rect 10 -23 17 -21
<< gv1 >>
rect -41 6 -36 11
rect -14 6 -9 11
rect 29 6 34 11
rect 17 -3 22 2
rect -41 -11 -36 -6
rect -14 -11 -9 -6
rect 29 -11 34 -6
rect -32 -22 -27 -17
rect 11 -22 16 -17
<< labels >>
rlabel gv1 -39 8 -38 9 1 Vdd!
rlabel polycontact -30 0 -29 1 1 a
rlabel metal1 -22 0 -21 1 1 na
rlabel gv1 -39 -9 -38 -8 1 GND!
rlabel polycontact 22 -21 23 -20 1 g1
rlabel polycontact -6 -27 -5 -26 1 g0
rlabel metal1 8 -1 9 0 1 out
<< end >>
