magic
tech scmos
timestamp 1757617612
<< pwell >>
rect -24 -13 12 3
<< nwell >>
rect -24 3 12 19
<< polysilicon >>
rect -5 15 0 17
rect -5 6 0 10
rect -5 -2 0 1
rect -5 -11 0 -7
<< ndiffusion >>
rect -13 -7 -12 -2
rect -7 -7 -5 -2
rect 0 -7 3 -2
rect 8 -7 9 -2
<< pdiffusion >>
rect -13 10 -12 15
rect -7 10 -5 15
rect 0 10 3 15
rect 8 10 9 15
<< metal1 >>
rect -17 10 -12 15
rect 3 -2 8 10
rect -17 -7 -12 -2
<< ntransistor >>
rect -5 -7 0 -2
<< ptransistor >>
rect -5 10 0 15
<< polycontact >>
rect -5 1 0 6
<< ndcontact >>
rect -12 -7 -7 -2
rect 3 -7 8 -2
<< pdcontact >>
rect -12 10 -7 15
rect 3 10 8 15
<< psubstratepcontact >>
rect -22 -7 -17 -2
<< nsubstratencontact >>
rect -22 10 -17 15
<< labels >>
rlabel polycontact -4 1 -3 2 1 in
rlabel nsubstratencontact -20 12 -19 13 3 Vdd!
rlabel psubstratepcontact -20 -5 -19 -4 3 GND!
rlabel metal1 6 2 7 3 7 out
<< end >>
