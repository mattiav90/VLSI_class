magic
tech scmos
timestamp 1759210043
<< nwell >>
rect -2 35 251 50
rect -1 24 251 35
rect -1 23 125 24
rect -1 20 124 23
rect 132 20 251 24
<< pwell >>
rect -1 11 124 20
rect 132 18 251 20
rect 131 16 251 18
rect -1 10 127 11
rect 129 10 251 16
rect -1 -3 251 10
<< metal1 >>
rect 66 46 161 49
rect 66 29 70 46
rect 106 36 113 43
rect 107 30 112 36
rect 24 15 27 20
rect 66 16 69 21
rect 108 17 111 22
rect 158 20 161 46
rect 195 21 197 23
rect 23 2 28 14
rect 125 6 127 11
rect 143 2 146 20
rect 194 18 211 21
rect 219 17 222 22
rect 23 -1 146 2
<< metal2 >>
rect 106 41 113 43
rect 106 38 247 41
rect 106 36 113 38
rect 6 28 12 33
rect 36 29 61 32
rect 79 29 104 32
rect 120 29 139 32
rect 175 28 207 31
rect 14 17 19 22
rect 31 16 38 23
rect 55 16 62 23
rect 73 16 80 23
rect 115 16 122 23
rect 243 19 247 38
rect 231 16 247 19
rect 7 10 13 11
rect 7 6 138 10
rect 176 9 208 12
<< gv1 >>
rect 107 37 112 42
<< metal3 >>
rect 34 34 103 37
rect 34 23 38 34
rect 100 23 103 34
rect 13 16 20 23
rect 31 16 38 23
rect 55 16 62 23
rect 73 16 80 23
rect 97 16 104 23
rect 115 16 122 23
rect 16 7 20 16
rect 55 7 59 16
rect 16 3 59 7
rect 76 7 80 16
rect 117 7 120 16
rect 76 3 120 7
<< gv2 >>
rect 14 17 19 22
rect 32 17 37 22
rect 56 17 61 22
rect 74 17 79 22
rect 98 17 103 22
rect 116 17 121 22
use nand2  nand2_3
timestamp 1759205441
transform 1 0 214 0 1 22
box -20 -22 30 16
use and2  and2_0
timestamp 1759209702
transform 1 0 147 0 1 22
box -21 -19 60 15
use nand2  nand2_0
timestamp 1759205441
transform 1 0 19 0 1 22
box -20 -22 30 16
use nand2  nand2_1
timestamp 1759205441
transform 1 0 61 0 1 22
box -20 -22 30 16
use nand2  nand2_2
timestamp 1759205441
transform 1 0 103 0 1 22
box -20 -22 30 16
<< labels >>
rlabel metal2 6 28 12 33 1 Vdd!
rlabel metal2 14 17 19 22 1 a
rlabel metal2 32 17 37 22 1 b
rlabel metal2 74 17 79 22 1 cin
rlabel metal1 24 15 27 20 1 ab
rlabel metal1 66 16 69 21 1 acin
rlabel metal1 108 17 111 22 1 bcin
rlabel metal2 10 7 13 11 1 GND!
rlabel metal1 195 18 197 23 1 andout
rlabel metal1 219 17 222 22 1 cout
<< end >>
