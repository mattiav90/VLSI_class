magic
tech scmos
timestamp 1759210717
use fuladdall  fuladdall_0
timestamp 1759210717
transform 1 0 3 0 1 2
box -3 -2 483 66
<< end >>
