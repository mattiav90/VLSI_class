magic
tech scmos
timestamp 1759205441
<< error_p >>
rect -12 10 24 11
rect 22 6 24 10
<< nwell >>
rect -20 -2 28 16
<< pwell >>
rect -20 -22 30 -2
<< ntransistor >>
rect -5 -16 0 -11
rect 13 -16 18 -11
<< ptransistor >>
rect -5 6 0 11
rect 13 6 18 11
<< ndiffusion >>
rect -7 -16 -5 -11
rect 0 -16 13 -11
rect 18 -16 19 -11
<< pdiffusion >>
rect -7 6 -5 11
rect 0 6 4 11
rect 9 6 13 11
rect 18 6 19 11
<< ndcontact >>
rect -12 -16 -7 -11
rect 19 -16 24 -11
<< pdcontact >>
rect -12 6 -7 11
rect 4 6 9 11
rect 19 6 24 11
<< polysilicon >>
rect -5 11 0 14
rect 13 11 18 14
rect -5 0 0 6
rect -5 -11 0 -5
rect 13 0 18 6
rect 13 -11 18 -5
rect -5 -19 0 -16
rect 13 -19 18 -16
<< polycontact >>
rect -5 -5 0 0
rect 13 -5 18 0
<< metal1 >>
rect -13 11 -6 12
rect 18 11 25 12
rect -13 6 -12 11
rect -7 6 -6 11
rect -13 5 -6 6
rect -6 0 1 1
rect -6 -5 -5 0
rect 0 -5 1 0
rect -6 -6 1 -5
rect -13 -11 -6 -10
rect -13 -16 -12 -11
rect -7 -16 -6 -11
rect 4 -11 9 6
rect 18 6 19 11
rect 24 6 25 11
rect 18 5 25 6
rect 12 0 19 1
rect 12 -5 13 0
rect 18 -5 19 0
rect 12 -6 19 -5
rect 4 -16 19 -11
rect -13 -17 -6 -16
<< metal2 >>
rect -13 10 -6 12
rect 18 10 25 12
rect -13 7 25 10
rect -13 5 -6 7
rect 18 5 25 7
rect -6 -6 1 1
rect 12 -6 19 1
rect -13 -17 -6 -10
<< gv1 >>
rect -12 6 -7 11
rect 19 6 24 11
rect -5 -5 0 0
rect 13 -5 18 0
rect -12 -16 -7 -11
<< labels >>
rlabel pdcontact -10 8 -9 9 1 Vdd!
rlabel polycontact -3 -3 -2 -2 1 a
rlabel gv1 -11 -14 -9 -13 1 GND!
rlabel metal1 6 -3 7 -2 1 out
rlabel polycontact 15 -3 16 -2 1 b
<< end >>
