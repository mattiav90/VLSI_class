magic
tech scmos
timestamp 1758854531
<< nwell >>
rect -2 31 264 57
<< pwell >>
rect -2 -2 264 31
<< ntransistor >>
rect 15 20 20 25
rect 40 20 44 25
rect 48 20 52 25
rect 59 20 63 25
rect 67 20 71 25
rect 102 20 107 25
rect 127 20 131 25
rect 135 20 139 25
rect 146 20 150 25
rect 154 20 158 25
rect 189 20 194 25
rect 214 20 218 25
rect 222 20 226 25
rect 233 20 237 25
rect 241 20 245 25
<< ptransistor >>
rect 15 37 20 42
rect 40 37 44 42
rect 48 37 52 42
rect 59 37 63 42
rect 67 37 71 42
rect 102 37 107 42
rect 127 37 131 42
rect 135 37 139 42
rect 146 37 150 42
rect 154 37 158 42
rect 189 37 194 42
rect 214 37 218 42
rect 222 37 226 42
rect 233 37 237 42
rect 241 37 245 42
<< ndiffusion >>
rect 11 20 15 25
rect 20 20 23 25
rect 32 20 33 25
rect 38 20 40 25
rect 44 20 48 25
rect 52 20 53 25
rect 58 20 59 25
rect 63 20 67 25
rect 71 20 76 25
rect 81 20 82 25
rect 98 20 102 25
rect 107 20 110 25
rect 119 20 120 25
rect 125 20 127 25
rect 131 20 135 25
rect 139 20 140 25
rect 145 20 146 25
rect 150 20 154 25
rect 158 20 163 25
rect 168 20 169 25
rect 185 20 189 25
rect 194 20 197 25
rect 206 20 207 25
rect 212 20 214 25
rect 218 20 222 25
rect 226 20 227 25
rect 232 20 233 25
rect 237 20 241 25
rect 245 20 250 25
rect 255 20 256 25
<< pdiffusion >>
rect 11 37 15 42
rect 20 37 23 42
rect 32 37 33 42
rect 38 37 40 42
rect 44 37 48 42
rect 52 37 53 42
rect 58 37 59 42
rect 63 37 67 42
rect 71 37 76 42
rect 81 37 82 42
rect 98 37 102 42
rect 107 37 110 42
rect 119 37 120 42
rect 125 37 127 42
rect 131 37 135 42
rect 139 37 140 42
rect 145 37 146 42
rect 150 37 154 42
rect 158 37 163 42
rect 168 37 169 42
rect 185 37 189 42
rect 194 37 197 42
rect 206 37 207 42
rect 212 37 214 42
rect 218 37 222 42
rect 226 37 227 42
rect 232 37 233 42
rect 237 37 241 42
rect 245 37 250 42
rect 255 37 256 42
<< ndcontact >>
rect 6 20 11 25
rect 23 20 28 25
rect 33 20 38 25
rect 53 20 58 25
rect 76 20 81 25
rect 93 20 98 25
rect 110 20 115 25
rect 120 20 125 25
rect 140 20 145 25
rect 163 20 168 25
rect 180 20 185 25
rect 197 20 202 25
rect 207 20 212 25
rect 227 20 232 25
rect 250 20 255 25
<< pdcontact >>
rect 6 37 11 42
rect 23 37 28 42
rect 33 37 38 42
rect 53 37 58 42
rect 76 37 81 42
rect 93 37 98 42
rect 110 37 115 42
rect 120 37 125 42
rect 140 37 145 42
rect 163 37 168 42
rect 180 37 185 42
rect 197 37 202 42
rect 207 37 212 42
rect 227 37 232 42
rect 250 37 255 42
<< polysilicon >>
rect 15 42 20 46
rect 40 42 44 47
rect 48 42 52 45
rect 59 42 63 45
rect 67 42 71 47
rect 102 42 107 46
rect 127 42 131 47
rect 135 42 139 45
rect 146 42 150 45
rect 154 42 158 47
rect 189 42 194 46
rect 214 42 218 47
rect 222 42 226 45
rect 233 42 237 45
rect 241 42 245 47
rect 15 34 20 37
rect 15 25 20 29
rect 40 25 44 37
rect 48 33 52 37
rect 59 33 63 37
rect 48 25 52 29
rect 59 25 63 29
rect 67 25 71 37
rect 102 34 107 37
rect 102 25 107 29
rect 127 25 131 37
rect 135 33 139 37
rect 146 33 150 37
rect 135 25 139 29
rect 146 25 150 29
rect 154 25 158 37
rect 189 34 194 37
rect 189 25 194 29
rect 214 25 218 37
rect 222 33 226 37
rect 233 33 237 37
rect 222 25 226 29
rect 233 25 237 29
rect 241 25 245 37
rect 15 14 20 20
rect 40 7 44 20
rect 48 17 52 20
rect 59 14 63 20
rect 67 13 71 20
rect 102 14 107 20
rect 127 7 131 20
rect 135 17 139 20
rect 146 14 150 20
rect 154 13 158 20
rect 189 14 194 20
rect 214 7 218 20
rect 222 17 226 20
rect 233 14 237 20
rect 241 13 245 20
<< polycontact >>
rect 48 45 53 50
rect 58 45 63 50
rect 135 45 140 50
rect 145 45 150 50
rect 222 45 227 50
rect 232 45 237 50
rect 15 29 20 34
rect 102 29 107 34
rect 189 29 194 34
rect 48 12 53 17
rect 58 9 63 14
rect 67 8 72 13
rect 135 12 140 17
rect 145 9 150 14
rect 154 8 159 13
rect 222 12 227 17
rect 232 9 237 14
rect 241 8 246 13
rect 39 2 44 7
rect 126 2 131 7
rect 213 2 218 7
<< metal1 >>
rect 50 54 111 57
rect 50 50 53 54
rect 17 47 48 50
rect 5 42 12 43
rect 5 37 6 42
rect 11 37 12 42
rect 5 36 12 37
rect 17 34 20 47
rect 58 50 88 51
rect 107 50 111 54
rect 145 50 175 51
rect 232 50 262 51
rect 63 48 88 50
rect 32 42 39 43
rect 75 42 82 43
rect 5 25 12 26
rect 5 20 6 25
rect 11 20 12 25
rect 5 19 12 20
rect 17 15 20 29
rect 25 25 28 37
rect 32 37 33 42
rect 38 37 39 42
rect 32 36 39 37
rect 54 31 58 37
rect 75 37 76 42
rect 81 37 82 42
rect 75 36 82 37
rect 63 31 70 34
rect 54 28 70 31
rect 25 16 28 20
rect 32 25 39 26
rect 54 25 58 28
rect 63 27 70 28
rect 32 20 33 25
rect 38 20 39 25
rect 75 25 82 26
rect 75 20 76 25
rect 81 20 82 25
rect 32 19 39 20
rect 75 19 82 20
rect 14 8 21 15
rect 25 13 48 16
rect 38 2 39 7
rect 50 3 53 12
rect 57 14 64 15
rect 57 9 58 14
rect 63 9 64 14
rect 57 8 64 9
rect 72 8 73 13
rect 85 3 88 48
rect 104 47 135 50
rect 92 42 99 43
rect 92 37 93 42
rect 98 37 99 42
rect 92 36 99 37
rect 104 34 107 47
rect 150 48 175 50
rect 119 42 126 43
rect 162 42 169 43
rect 92 25 99 26
rect 92 20 93 25
rect 98 20 99 25
rect 92 19 99 20
rect 104 15 107 29
rect 112 25 115 37
rect 119 37 120 42
rect 125 37 126 42
rect 119 36 126 37
rect 141 31 145 37
rect 162 37 163 42
rect 168 37 169 42
rect 162 36 169 37
rect 150 31 157 34
rect 141 28 157 31
rect 112 16 115 20
rect 119 25 126 26
rect 141 25 145 28
rect 150 27 157 28
rect 119 20 120 25
rect 125 20 126 25
rect 162 25 169 26
rect 162 20 163 25
rect 168 20 169 25
rect 119 19 126 20
rect 162 19 169 20
rect 101 8 108 15
rect 112 13 135 16
rect 50 0 88 3
rect 125 2 126 7
rect 137 3 140 12
rect 144 14 151 15
rect 144 9 145 14
rect 150 9 151 14
rect 144 8 151 9
rect 159 8 160 13
rect 172 3 175 48
rect 191 47 222 50
rect 179 42 186 43
rect 179 37 180 42
rect 185 37 186 42
rect 179 36 186 37
rect 191 34 194 47
rect 237 48 262 50
rect 206 42 213 43
rect 249 42 256 43
rect 179 25 186 26
rect 179 20 180 25
rect 185 20 186 25
rect 179 19 186 20
rect 191 15 194 29
rect 199 25 202 37
rect 206 37 207 42
rect 212 37 213 42
rect 206 36 213 37
rect 228 31 232 37
rect 249 37 250 42
rect 255 37 256 42
rect 249 36 256 37
rect 237 31 244 34
rect 228 28 244 31
rect 199 16 202 20
rect 206 25 213 26
rect 228 25 232 28
rect 237 27 244 28
rect 206 20 207 25
rect 212 20 213 25
rect 249 25 256 26
rect 249 20 250 25
rect 255 20 256 25
rect 206 19 213 20
rect 249 19 256 20
rect 188 8 195 15
rect 199 13 222 16
rect 137 0 175 3
rect 212 2 213 7
rect 218 2 219 6
rect 212 -1 219 2
rect 224 3 227 12
rect 231 14 238 15
rect 231 9 232 14
rect 237 9 238 14
rect 242 13 250 15
rect 231 8 238 9
rect 246 8 250 13
rect 242 7 250 8
rect 259 3 262 48
rect 224 0 262 3
<< metal2 >>
rect -2 42 1 57
rect 5 42 12 43
rect 32 42 39 43
rect 75 42 82 43
rect 92 42 99 43
rect 119 42 126 43
rect 162 42 169 43
rect 179 42 186 43
rect 206 42 213 43
rect 249 42 256 43
rect -2 38 256 42
rect -2 37 58 38
rect -2 -2 1 37
rect 5 36 12 37
rect 32 36 39 37
rect 75 36 82 38
rect 92 37 145 38
rect 162 37 232 38
rect 92 36 99 37
rect 119 36 126 37
rect 162 36 169 37
rect 179 36 186 37
rect 206 36 213 37
rect 249 36 256 38
rect 63 27 70 34
rect 150 27 157 34
rect 237 27 244 34
rect 5 25 12 26
rect 32 25 39 26
rect 5 23 58 25
rect 75 24 82 26
rect 92 25 99 26
rect 119 25 126 26
rect 92 24 145 25
rect 75 23 145 24
rect 162 24 169 26
rect 179 25 186 26
rect 206 25 213 26
rect 179 24 232 25
rect 162 23 232 24
rect 249 23 256 26
rect 260 23 263 57
rect 5 20 263 23
rect 5 19 12 20
rect 32 19 39 20
rect 75 19 82 20
rect 92 19 99 20
rect 119 19 126 20
rect 162 19 169 20
rect 179 19 186 20
rect 206 19 213 20
rect 249 19 256 20
rect 14 14 21 15
rect 57 14 64 15
rect 14 10 64 14
rect 14 8 21 10
rect 57 8 64 10
rect 101 14 108 15
rect 144 14 151 15
rect 101 10 151 14
rect 101 8 108 10
rect 144 8 151 10
rect 188 14 195 15
rect 231 14 238 15
rect 188 10 238 14
rect 188 8 195 10
rect 231 8 238 10
rect 242 7 250 15
rect 212 -1 219 6
rect 260 -2 263 20
<< gv1 >>
rect 6 37 11 42
rect 33 37 38 42
rect 76 37 81 42
rect 93 37 98 42
rect 120 37 125 42
rect 163 37 168 42
rect 180 37 185 42
rect 207 37 212 42
rect 250 37 255 42
rect 64 28 69 33
rect 151 28 156 33
rect 238 28 243 33
rect 6 20 11 25
rect 33 20 38 25
rect 76 20 81 25
rect 93 20 98 25
rect 120 20 125 25
rect 163 20 168 25
rect 180 20 185 25
rect 207 20 212 25
rect 250 20 255 25
rect 15 9 20 14
rect 58 9 63 14
rect 102 9 107 14
rect 145 9 150 14
rect 189 9 194 14
rect 232 9 237 14
rect 243 8 249 14
rect 213 0 218 5
<< metal3 >>
rect 63 27 70 34
rect 150 32 157 34
rect 150 28 226 32
rect 150 27 157 28
rect 64 4 69 27
rect 223 12 226 28
rect 242 12 250 15
rect 223 9 250 12
rect 242 7 250 9
rect 212 4 219 6
rect 64 0 219 4
rect 212 -1 219 0
<< gv2 >>
rect 64 28 69 33
rect 151 28 156 33
rect 243 8 249 14
rect 213 0 218 5
<< labels >>
rlabel metal1 41 4 42 5 1 g0
rlabel polycontact 41 4 42 5 1 2lut_0/g0
rlabel gv2 66 30 67 31 1 out0
rlabel metal1 191 31 192 32 1 a
rlabel metal1 69 10 70 11 1 g1
rlabel metal1 156 10 157 11 1 g3
rlabel metal1 229 30 230 31 1 out
rlabel polycontact 191 31 192 32 1 2lut_2/a
rlabel metal1 199 31 200 32 1 2lut_2/na
rlabel gv1 182 22 183 23 1 2lut_2/GND!
rlabel metal1 229 30 230 31 1 2lut_2/out
rlabel polycontact 104 31 105 32 1 2lut_1/a
rlabel metal1 112 31 113 32 1 2lut_1/na
rlabel gv1 95 22 96 23 1 2lut_1/GND!
rlabel polycontact 156 10 157 11 1 2lut_1/g1
rlabel polycontact 69 10 70 11 1 2lut_0/g1
rlabel metal1 55 30 56 31 1 2lut_0/out
rlabel metal1 142 30 143 31 1 2lut_1/out
rlabel gv2 153 30 154 31 1 out1
rlabel gv1 8 22 9 23 1 2lut_0/GND!
rlabel metal1 25 31 26 32 1 2lut_0/na
rlabel polycontact 17 31 18 32 1 2lut_0/a
rlabel polycontact 128 4 129 5 1 2lut_1/g0
rlabel gv1 95 39 96 40 1 2lut_1/Vdd!
rlabel polycontact 215 4 216 5 1 2lut_2/g0
rlabel polycontact 243 10 244 11 1 2lut_2/g1
rlabel gv1 182 39 183 40 1 2lut_2/Vdd!
rlabel metal1 128 4 129 5 1 g2
rlabel metal1 17 31 18 32 1 b
rlabel metal2 8 22 9 23 1 GND!
rlabel gv1 8 39 9 40 1 2lut_0/Vdd!
rlabel metal2 8 39 9 40 1 Vdd!
<< end >>
