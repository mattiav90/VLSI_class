magic
tech scmos
timestamp 1757627839
<< nwell >>
rect -24 -2 28 15
<< pwell >>
rect -24 -19 28 -2
<< ntransistor >>
rect -5 -13 0 -8
rect 11 -13 16 -8
<< ptransistor >>
rect -5 4 0 9
rect 11 4 16 9
<< ndiffusion >>
rect -7 -13 -5 -8
rect 0 -13 11 -8
rect 16 -13 17 -8
<< pdiffusion >>
rect -7 4 -5 9
rect 0 4 3 9
rect 8 4 11 9
rect 16 4 17 9
<< ndcontact >>
rect -12 -13 -7 -8
rect 17 -13 22 -8
<< pdcontact >>
rect -12 4 -7 9
rect 3 4 8 9
rect 17 4 22 9
<< psubstratepcontact >>
rect -21 -13 -16 -8
<< nsubstratencontact >>
rect -21 4 -16 9
<< polysilicon >>
rect -5 9 0 12
rect 11 9 16 12
rect -5 0 0 4
rect -5 -8 0 -5
rect 11 0 16 4
rect 11 -8 16 -5
rect -5 -16 0 -13
rect 11 -16 16 -13
<< polycontact >>
rect -5 -5 0 0
rect 11 -5 16 0
<< metal1 >>
rect -12 12 22 15
rect -12 9 -7 12
rect 17 9 22 12
rect -16 4 -12 9
rect 3 -8 8 4
rect -16 -13 -12 -8
rect 3 -13 17 -8
<< labels >>
rlabel metal1 5 -3 6 -2 1 out
rlabel pdcontact -10 6 -9 7 1 Vdd!
rlabel psubstratepcontact -19 -11 -18 -10 1 GND!
rlabel polycontact -3 -3 -2 -2 1 a
rlabel polycontact 13 -3 14 -2 1 b
<< end >>
