magic
tech scmos
timestamp 1760051112
<< pwell >>
rect 99 15 107 17
rect 107 10 112 11
rect 101 8 112 10
rect 101 0 122 8
rect 224 0 233 6
<< metal2 >>
rect -5 45 2 52
rect 97 46 132 49
rect 4 34 11 41
rect 90 34 97 41
rect 167 31 174 38
rect -5 21 2 28
rect 96 24 131 27
<< metal3 >>
rect 4 34 11 41
rect 45 31 52 38
rect 90 34 97 41
rect 212 34 219 41
rect 100 11 107 15
rect 100 8 134 11
<< gv2 >>
rect 46 32 51 37
<< metal4 >>
rect 45 31 52 38
rect 48 17 52 31
rect 48 13 107 17
rect 100 8 107 13
<< gv3 >>
rect 46 32 51 37
rect 101 9 106 14
use xor2  xor2_0
timestamp 1759199526
transform 1 0 30 0 1 44
box -41 -44 81 23
use xor2  xor2_1
timestamp 1759199526
transform 1 0 152 0 1 44
box -41 -44 81 23
<< labels >>
rlabel metal3 7 37 8 38 1 a
rlabel metal3 93 37 94 38 1 b
rlabel metal3 215 37 216 38 1 cin
rlabel metal2 170 34 171 35 1 out
rlabel metal2 -2 48 -1 49 1 Vdd!
rlabel metal2 -2 24 -1 25 1 GND!
rlabel gv2 47 33 49 35 1 mid
<< end >>
