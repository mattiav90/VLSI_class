magic
tech scmos
timestamp 1760053292
<< nwell >>
rect -247 39 7 47
<< pwell >>
rect -10 -21 249 -1
<< metal1 >>
rect 218 9 221 14
<< metal2 >>
rect -239 26 -235 30
rect -18 25 9 29
rect -68 11 -63 16
rect -239 2 -236 5
rect -16 3 9 6
<< metal3 >>
rect -230 14 -227 19
rect -23 14 -18 19
rect 71 13 78 20
rect -207 -17 -203 -10
rect 14 -17 17 3
rect -207 -20 17 -17
<< metal4 >>
rect -142 42 33 45
rect -142 20 -139 42
rect 30 20 33 42
rect -146 13 -139 20
rect -24 13 -17 20
rect 29 13 36 20
rect 71 13 78 20
rect -21 -13 -17 13
rect 73 -13 76 13
rect -21 -16 76 -13
<< gv3 >>
rect -145 14 -140 19
rect -23 14 -18 19
rect 30 14 35 19
rect 72 14 77 19
use sum  sum_0
timestamp 1760051112
transform 1 0 -236 0 1 -21
box -11 0 233 67
use cout  cout_0
timestamp 1760046497
transform 1 0 -2 0 1 -3
box -2 -3 251 50
<< labels >>
rlabel metal3 -229 16 -228 17 1 a
rlabel gv3 -143 16 -142 17 1 b
rlabel gv3 -21 16 -20 17 1 cin
rlabel space -247 -21 -125 46 1 Vdd!
rlabel metal2 -238 3 -237 4 1 GND!
rlabel metal2 -66 13 -65 15 1 sum
rlabel metal1 218 11 219 12 1 cout
rlabel metal2 -238 27 -237 28 1 Vdd!
<< end >>
