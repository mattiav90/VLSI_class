magic
tech scmos
timestamp 1757968460
<< nwell >>
rect -17 17 332 20
rect -17 15 281 17
rect -17 2 80 15
rect 132 2 229 15
rect 317 8 321 17
<< pwell >>
rect -17 -13 80 2
rect 83 -13 88 -4
rect 132 -12 229 2
rect 101 -13 229 -12
rect 232 -13 237 -4
rect 250 -13 281 -12
rect -17 -16 289 -13
<< ntransistor >>
rect -5 -9 0 -4
rect 11 -9 16 -4
rect 43 -9 48 -4
rect 59 -9 64 -4
rect 144 -9 149 -4
rect 160 -9 165 -4
rect 192 -9 197 -4
rect 208 -9 213 -4
<< ptransistor >>
rect -5 8 0 13
rect 11 8 16 13
rect 43 8 48 13
rect 59 8 64 13
rect 144 8 149 13
rect 160 8 165 13
rect 192 8 197 13
rect 208 8 213 13
<< ndiffusion >>
rect -6 -9 -5 -4
rect 0 -9 3 -4
rect 8 -9 11 -4
rect 16 -9 17 -4
rect 42 -9 43 -4
rect 48 -9 51 -4
rect 56 -9 59 -4
rect 64 -9 65 -4
rect 143 -9 144 -4
rect 149 -9 152 -4
rect 157 -9 160 -4
rect 165 -9 166 -4
rect 191 -9 192 -4
rect 197 -9 200 -4
rect 205 -9 208 -4
rect 213 -9 214 -4
<< pdiffusion >>
rect -6 8 -5 13
rect 0 8 11 13
rect 16 8 17 13
rect 42 8 43 13
rect 48 8 59 13
rect 64 8 65 13
rect 143 8 144 13
rect 149 8 160 13
rect 165 8 166 13
rect 191 8 192 13
rect 197 8 208 13
rect 213 8 214 13
<< ndcontact >>
rect -11 -9 -6 -4
rect 3 -9 8 -4
rect 17 -9 22 -4
rect 37 -9 42 -4
rect 51 -9 56 -4
rect 65 -9 70 -4
rect 138 -9 143 -4
rect 152 -9 157 -4
rect 166 -9 171 -4
rect 186 -9 191 -4
rect 200 -9 205 -4
rect 214 -9 219 -4
<< pdcontact >>
rect -11 8 -6 13
rect 17 8 22 13
rect 37 8 42 13
rect 65 8 70 13
rect 138 8 143 13
rect 166 8 171 13
rect 186 8 191 13
rect 214 8 219 13
<< psubstratepcontact >>
rect 26 -9 31 -4
rect 74 -9 79 -4
rect 175 -9 180 -4
rect 223 -9 228 -4
<< nsubstratencontact >>
rect 26 8 31 13
rect 74 8 79 13
rect 175 8 180 13
rect 223 8 228 13
<< polysilicon >>
rect -5 13 0 17
rect 11 13 16 17
rect 43 13 48 17
rect 59 13 64 17
rect 144 13 149 17
rect 160 13 165 17
rect 192 13 197 17
rect 208 13 213 17
rect -5 4 0 8
rect -5 -4 0 -1
rect 11 4 16 8
rect 11 -4 16 -1
rect 43 4 48 8
rect 43 -4 48 -1
rect 59 4 64 8
rect 59 -4 64 -1
rect 144 4 149 8
rect 144 -4 149 -1
rect 160 4 165 8
rect 160 -4 165 -1
rect 192 4 197 8
rect 192 -4 197 -1
rect 208 4 213 8
rect 208 -4 213 -1
rect -5 -12 0 -9
rect 11 -12 16 -9
rect 43 -12 48 -9
rect 59 -12 64 -9
rect 144 -12 149 -9
rect 160 -12 165 -9
rect 192 -12 197 -9
rect 208 -12 213 -9
<< polycontact >>
rect -5 -1 0 4
rect 11 -1 16 4
rect 43 -1 48 4
rect 59 -1 64 4
rect 144 -1 149 4
rect 160 -1 165 4
rect 192 -1 197 4
rect 208 -1 213 4
<< metal1 >>
rect 26 17 321 20
rect 26 16 96 17
rect 175 16 245 17
rect 26 13 31 16
rect 74 13 79 16
rect 175 13 180 16
rect 223 13 228 16
rect -6 8 8 13
rect 22 8 26 13
rect 42 8 51 13
rect 70 8 74 13
rect 143 8 157 13
rect 171 8 175 13
rect 191 8 200 13
rect 219 8 223 13
rect 317 8 321 17
rect 3 4 8 8
rect 11 4 16 5
rect 43 4 48 5
rect 3 -4 8 -1
rect 51 -4 56 8
rect 59 4 64 5
rect 152 4 157 8
rect 160 4 165 5
rect 192 4 197 5
rect 152 -4 157 -1
rect 200 -4 205 8
rect 208 4 213 5
rect 292 -1 298 4
rect 302 0 305 3
rect 309 -1 315 4
rect 22 -9 26 -4
rect 70 -9 74 -4
rect -11 -13 -6 -9
rect 17 -13 22 -9
rect 37 -13 42 -9
rect 65 -13 70 -9
rect 83 -13 88 -4
rect 171 -9 175 -4
rect 219 -9 223 -4
rect 138 -13 143 -9
rect 166 -13 171 -9
rect 186 -13 191 -9
rect 214 -13 219 -9
rect 232 -13 237 -4
rect -11 -16 289 -13
<< m2contact >>
rect 51 8 56 13
rect 200 8 205 13
rect 3 -1 8 4
rect 94 -1 99 4
rect 107 -1 112 4
rect 120 -1 125 4
rect 152 -1 157 4
rect 243 -1 248 4
rect 256 -1 261 4
rect 269 -1 274 4
rect 287 -1 292 4
rect 315 -1 320 4
<< metal2 >>
rect 56 8 125 13
rect 205 8 274 13
rect 120 4 125 8
rect 269 4 274 8
rect 8 -1 94 4
rect 157 -1 243 4
rect 107 -12 112 -1
rect 256 -5 261 -1
rect 287 -5 292 -1
rect 256 -8 292 -5
rect 315 -12 320 -1
rect 107 -16 320 -12
use nor2  nor2_0 ../nor2
timestamp 1757643574
transform 1 0 298 0 1 4
box -17 -20 34 15
use nand2  nand2_1 ../nand2
timestamp 1757633819
transform 1 0 253 0 1 4
box -24 -19 28 15
use nand2  nand2_0
timestamp 1757633819
transform 1 0 104 0 1 4
box -24 -19 28 15
<< labels >>
rlabel polycontact -4 1 -3 2 1 in1
rlabel metal1 12 4 13 5 1 in2
rlabel metal1 45 4 46 5 1 in3
rlabel metal1 62 4 63 5 1 in4
rlabel polycontact 146 1 146 2 1 in5
rlabel metal1 162 4 163 5 1 in6
rlabel metal1 193 4 194 5 1 in7
rlabel metal1 209 4 210 5 1 in8
rlabel metal1 19 -15 21 -14 1 GND!
rlabel metal1 43 -15 44 -14 1 GND!
rlabel m2contact 109 1 110 3 1 out4_1
rlabel m2contact 257 1 259 2 1 out4_2
rlabel metal1 303 1 304 3 1 out
<< end >>
