magic
tech scmos
timestamp 1759210420
<< pwell >>
rect 223 15 317 36
rect 223 -2 483 15
<< metal2 >>
rect 4 44 10 49
rect 102 44 126 47
rect 218 44 242 47
rect 169 30 173 35
rect 4 20 9 25
rect 105 22 129 25
rect 222 22 246 25
<< metal3 >>
rect 13 33 18 38
rect 53 29 60 36
rect 99 33 104 38
rect 126 32 133 39
rect 213 33 218 38
<< gv2 >>
rect 54 30 59 35
rect 127 33 132 38
<< metal4 >>
rect 53 29 60 36
rect 57 16 60 29
rect 126 32 133 39
rect 126 16 129 32
rect 57 13 129 16
<< gv3 >>
rect 54 30 59 35
rect 127 33 132 38
use cout  cout_0
timestamp 1759210420
transform 1 0 232 0 1 16
box -2 -3 251 50
use xor2  xor2_1
timestamp 1759199526
transform 1 0 152 0 1 42
box -41 -44 81 23
use xor2  xor2_0
timestamp 1759199526
transform 1 0 38 0 1 42
box -41 -44 81 23
<< labels >>
rlabel metal3 14 33 16 36 1 a
rlabel metal3 100 34 102 37 1 b
rlabel metal3 215 34 217 37 1 cin
rlabel metal2 169 30 173 35 1 out
rlabel metal2 4 44 10 49 1 Vdd!
rlabel metal2 4 20 9 25 1 GND!
<< end >>
