magic
tech scmos
timestamp 1758863309
<< nwell >>
rect -2 444 263 470
rect -2 385 263 411
rect -2 326 263 352
rect -2 267 263 293
rect -2 208 263 234
rect -2 149 263 175
rect -2 90 263 116
rect -2 31 263 57
<< pwell >>
rect -2 411 263 444
rect -2 352 263 385
rect -2 293 263 326
rect -2 234 263 267
rect -2 175 263 208
rect -2 116 263 149
rect -2 57 263 90
rect -2 -2 263 31
<< ntransistor >>
rect 15 433 20 438
rect 40 433 44 438
rect 48 433 52 438
rect 59 433 63 438
rect 67 433 71 438
rect 102 433 107 438
rect 127 433 131 438
rect 135 433 139 438
rect 146 433 150 438
rect 154 433 158 438
rect 189 433 194 438
rect 214 433 218 438
rect 222 433 226 438
rect 233 433 237 438
rect 241 433 245 438
rect 15 374 20 379
rect 40 374 44 379
rect 48 374 52 379
rect 59 374 63 379
rect 67 374 71 379
rect 102 374 107 379
rect 127 374 131 379
rect 135 374 139 379
rect 146 374 150 379
rect 154 374 158 379
rect 189 374 194 379
rect 214 374 218 379
rect 222 374 226 379
rect 233 374 237 379
rect 241 374 245 379
rect 15 315 20 320
rect 40 315 44 320
rect 48 315 52 320
rect 59 315 63 320
rect 67 315 71 320
rect 102 315 107 320
rect 127 315 131 320
rect 135 315 139 320
rect 146 315 150 320
rect 154 315 158 320
rect 189 315 194 320
rect 214 315 218 320
rect 222 315 226 320
rect 233 315 237 320
rect 241 315 245 320
rect 15 256 20 261
rect 40 256 44 261
rect 48 256 52 261
rect 59 256 63 261
rect 67 256 71 261
rect 102 256 107 261
rect 127 256 131 261
rect 135 256 139 261
rect 146 256 150 261
rect 154 256 158 261
rect 189 256 194 261
rect 214 256 218 261
rect 222 256 226 261
rect 233 256 237 261
rect 241 256 245 261
rect 15 197 20 202
rect 40 197 44 202
rect 48 197 52 202
rect 59 197 63 202
rect 67 197 71 202
rect 102 197 107 202
rect 127 197 131 202
rect 135 197 139 202
rect 146 197 150 202
rect 154 197 158 202
rect 189 197 194 202
rect 214 197 218 202
rect 222 197 226 202
rect 233 197 237 202
rect 241 197 245 202
rect 15 138 20 143
rect 40 138 44 143
rect 48 138 52 143
rect 59 138 63 143
rect 67 138 71 143
rect 102 138 107 143
rect 127 138 131 143
rect 135 138 139 143
rect 146 138 150 143
rect 154 138 158 143
rect 189 138 194 143
rect 214 138 218 143
rect 222 138 226 143
rect 233 138 237 143
rect 241 138 245 143
rect 15 79 20 84
rect 40 79 44 84
rect 48 79 52 84
rect 59 79 63 84
rect 67 79 71 84
rect 102 79 107 84
rect 127 79 131 84
rect 135 79 139 84
rect 146 79 150 84
rect 154 79 158 84
rect 189 79 194 84
rect 214 79 218 84
rect 222 79 226 84
rect 233 79 237 84
rect 241 79 245 84
rect 15 20 20 25
rect 40 20 44 25
rect 48 20 52 25
rect 59 20 63 25
rect 67 20 71 25
rect 102 20 107 25
rect 127 20 131 25
rect 135 20 139 25
rect 146 20 150 25
rect 154 20 158 25
rect 189 20 194 25
rect 214 20 218 25
rect 222 20 226 25
rect 233 20 237 25
rect 241 20 245 25
<< ptransistor >>
rect 15 450 20 455
rect 40 450 44 455
rect 48 450 52 455
rect 59 450 63 455
rect 67 450 71 455
rect 102 450 107 455
rect 127 450 131 455
rect 135 450 139 455
rect 146 450 150 455
rect 154 450 158 455
rect 189 450 194 455
rect 214 450 218 455
rect 222 450 226 455
rect 233 450 237 455
rect 241 450 245 455
rect 15 391 20 396
rect 40 391 44 396
rect 48 391 52 396
rect 59 391 63 396
rect 67 391 71 396
rect 102 391 107 396
rect 127 391 131 396
rect 135 391 139 396
rect 146 391 150 396
rect 154 391 158 396
rect 189 391 194 396
rect 214 391 218 396
rect 222 391 226 396
rect 233 391 237 396
rect 241 391 245 396
rect 15 332 20 337
rect 40 332 44 337
rect 48 332 52 337
rect 59 332 63 337
rect 67 332 71 337
rect 102 332 107 337
rect 127 332 131 337
rect 135 332 139 337
rect 146 332 150 337
rect 154 332 158 337
rect 189 332 194 337
rect 214 332 218 337
rect 222 332 226 337
rect 233 332 237 337
rect 241 332 245 337
rect 15 273 20 278
rect 40 273 44 278
rect 48 273 52 278
rect 59 273 63 278
rect 67 273 71 278
rect 102 273 107 278
rect 127 273 131 278
rect 135 273 139 278
rect 146 273 150 278
rect 154 273 158 278
rect 189 273 194 278
rect 214 273 218 278
rect 222 273 226 278
rect 233 273 237 278
rect 241 273 245 278
rect 15 214 20 219
rect 40 214 44 219
rect 48 214 52 219
rect 59 214 63 219
rect 67 214 71 219
rect 102 214 107 219
rect 127 214 131 219
rect 135 214 139 219
rect 146 214 150 219
rect 154 214 158 219
rect 189 214 194 219
rect 214 214 218 219
rect 222 214 226 219
rect 233 214 237 219
rect 241 214 245 219
rect 15 155 20 160
rect 40 155 44 160
rect 48 155 52 160
rect 59 155 63 160
rect 67 155 71 160
rect 102 155 107 160
rect 127 155 131 160
rect 135 155 139 160
rect 146 155 150 160
rect 154 155 158 160
rect 189 155 194 160
rect 214 155 218 160
rect 222 155 226 160
rect 233 155 237 160
rect 241 155 245 160
rect 15 96 20 101
rect 40 96 44 101
rect 48 96 52 101
rect 59 96 63 101
rect 67 96 71 101
rect 102 96 107 101
rect 127 96 131 101
rect 135 96 139 101
rect 146 96 150 101
rect 154 96 158 101
rect 189 96 194 101
rect 214 96 218 101
rect 222 96 226 101
rect 233 96 237 101
rect 241 96 245 101
rect 15 37 20 42
rect 40 37 44 42
rect 48 37 52 42
rect 59 37 63 42
rect 67 37 71 42
rect 102 37 107 42
rect 127 37 131 42
rect 135 37 139 42
rect 146 37 150 42
rect 154 37 158 42
rect 189 37 194 42
rect 214 37 218 42
rect 222 37 226 42
rect 233 37 237 42
rect 241 37 245 42
<< ndiffusion >>
rect 11 433 15 438
rect 20 433 23 438
rect 32 433 33 438
rect 38 433 40 438
rect 44 433 48 438
rect 52 433 53 438
rect 58 433 59 438
rect 63 433 67 438
rect 71 433 76 438
rect 81 433 82 438
rect 98 433 102 438
rect 107 433 110 438
rect 119 433 120 438
rect 125 433 127 438
rect 131 433 135 438
rect 139 433 140 438
rect 145 433 146 438
rect 150 433 154 438
rect 158 433 163 438
rect 168 433 169 438
rect 185 433 189 438
rect 194 433 197 438
rect 206 433 207 438
rect 212 433 214 438
rect 218 433 222 438
rect 226 433 227 438
rect 232 433 233 438
rect 237 433 241 438
rect 245 433 250 438
rect 255 433 256 438
rect 11 374 15 379
rect 20 374 23 379
rect 32 374 33 379
rect 38 374 40 379
rect 44 374 48 379
rect 52 374 53 379
rect 58 374 59 379
rect 63 374 67 379
rect 71 374 76 379
rect 81 374 82 379
rect 98 374 102 379
rect 107 374 110 379
rect 119 374 120 379
rect 125 374 127 379
rect 131 374 135 379
rect 139 374 140 379
rect 145 374 146 379
rect 150 374 154 379
rect 158 374 163 379
rect 168 374 169 379
rect 185 374 189 379
rect 194 374 197 379
rect 206 374 207 379
rect 212 374 214 379
rect 218 374 222 379
rect 226 374 227 379
rect 232 374 233 379
rect 237 374 241 379
rect 245 374 250 379
rect 255 374 256 379
rect 11 315 15 320
rect 20 315 23 320
rect 32 315 33 320
rect 38 315 40 320
rect 44 315 48 320
rect 52 315 53 320
rect 58 315 59 320
rect 63 315 67 320
rect 71 315 76 320
rect 81 315 82 320
rect 98 315 102 320
rect 107 315 110 320
rect 119 315 120 320
rect 125 315 127 320
rect 131 315 135 320
rect 139 315 140 320
rect 145 315 146 320
rect 150 315 154 320
rect 158 315 163 320
rect 168 315 169 320
rect 185 315 189 320
rect 194 315 197 320
rect 206 315 207 320
rect 212 315 214 320
rect 218 315 222 320
rect 226 315 227 320
rect 232 315 233 320
rect 237 315 241 320
rect 245 315 250 320
rect 255 315 256 320
rect 11 256 15 261
rect 20 256 23 261
rect 32 256 33 261
rect 38 256 40 261
rect 44 256 48 261
rect 52 256 53 261
rect 58 256 59 261
rect 63 256 67 261
rect 71 256 76 261
rect 81 256 82 261
rect 98 256 102 261
rect 107 256 110 261
rect 119 256 120 261
rect 125 256 127 261
rect 131 256 135 261
rect 139 256 140 261
rect 145 256 146 261
rect 150 256 154 261
rect 158 256 163 261
rect 168 256 169 261
rect 185 256 189 261
rect 194 256 197 261
rect 206 256 207 261
rect 212 256 214 261
rect 218 256 222 261
rect 226 256 227 261
rect 232 256 233 261
rect 237 256 241 261
rect 245 256 250 261
rect 255 256 256 261
rect 11 197 15 202
rect 20 197 23 202
rect 32 197 33 202
rect 38 197 40 202
rect 44 197 48 202
rect 52 197 53 202
rect 58 197 59 202
rect 63 197 67 202
rect 71 197 76 202
rect 81 197 82 202
rect 98 197 102 202
rect 107 197 110 202
rect 119 197 120 202
rect 125 197 127 202
rect 131 197 135 202
rect 139 197 140 202
rect 145 197 146 202
rect 150 197 154 202
rect 158 197 163 202
rect 168 197 169 202
rect 185 197 189 202
rect 194 197 197 202
rect 206 197 207 202
rect 212 197 214 202
rect 218 197 222 202
rect 226 197 227 202
rect 232 197 233 202
rect 237 197 241 202
rect 245 197 250 202
rect 255 197 256 202
rect 11 138 15 143
rect 20 138 23 143
rect 32 138 33 143
rect 38 138 40 143
rect 44 138 48 143
rect 52 138 53 143
rect 58 138 59 143
rect 63 138 67 143
rect 71 138 76 143
rect 81 138 82 143
rect 98 138 102 143
rect 107 138 110 143
rect 119 138 120 143
rect 125 138 127 143
rect 131 138 135 143
rect 139 138 140 143
rect 145 138 146 143
rect 150 138 154 143
rect 158 138 163 143
rect 168 138 169 143
rect 185 138 189 143
rect 194 138 197 143
rect 206 138 207 143
rect 212 138 214 143
rect 218 138 222 143
rect 226 138 227 143
rect 232 138 233 143
rect 237 138 241 143
rect 245 138 250 143
rect 255 138 256 143
rect 11 79 15 84
rect 20 79 23 84
rect 32 79 33 84
rect 38 79 40 84
rect 44 79 48 84
rect 52 79 53 84
rect 58 79 59 84
rect 63 79 67 84
rect 71 79 76 84
rect 81 79 82 84
rect 98 79 102 84
rect 107 79 110 84
rect 119 79 120 84
rect 125 79 127 84
rect 131 79 135 84
rect 139 79 140 84
rect 145 79 146 84
rect 150 79 154 84
rect 158 79 163 84
rect 168 79 169 84
rect 185 79 189 84
rect 194 79 197 84
rect 206 79 207 84
rect 212 79 214 84
rect 218 79 222 84
rect 226 79 227 84
rect 232 79 233 84
rect 237 79 241 84
rect 245 79 250 84
rect 255 79 256 84
rect 11 20 15 25
rect 20 20 23 25
rect 32 20 33 25
rect 38 20 40 25
rect 44 20 48 25
rect 52 20 53 25
rect 58 20 59 25
rect 63 20 67 25
rect 71 20 76 25
rect 81 20 82 25
rect 98 20 102 25
rect 107 20 110 25
rect 119 20 120 25
rect 125 20 127 25
rect 131 20 135 25
rect 139 20 140 25
rect 145 20 146 25
rect 150 20 154 25
rect 158 20 163 25
rect 168 20 169 25
rect 185 20 189 25
rect 194 20 197 25
rect 206 20 207 25
rect 212 20 214 25
rect 218 20 222 25
rect 226 20 227 25
rect 232 20 233 25
rect 237 20 241 25
rect 245 20 250 25
rect 255 20 256 25
<< pdiffusion >>
rect 11 450 15 455
rect 20 450 23 455
rect 32 450 33 455
rect 38 450 40 455
rect 44 450 48 455
rect 52 450 53 455
rect 58 450 59 455
rect 63 450 67 455
rect 71 450 76 455
rect 81 450 82 455
rect 98 450 102 455
rect 107 450 110 455
rect 119 450 120 455
rect 125 450 127 455
rect 131 450 135 455
rect 139 450 140 455
rect 145 450 146 455
rect 150 450 154 455
rect 158 450 163 455
rect 168 450 169 455
rect 185 450 189 455
rect 194 450 197 455
rect 206 450 207 455
rect 212 450 214 455
rect 218 450 222 455
rect 226 450 227 455
rect 232 450 233 455
rect 237 450 241 455
rect 245 450 250 455
rect 255 450 256 455
rect 11 391 15 396
rect 20 391 23 396
rect 32 391 33 396
rect 38 391 40 396
rect 44 391 48 396
rect 52 391 53 396
rect 58 391 59 396
rect 63 391 67 396
rect 71 391 76 396
rect 81 391 82 396
rect 98 391 102 396
rect 107 391 110 396
rect 119 391 120 396
rect 125 391 127 396
rect 131 391 135 396
rect 139 391 140 396
rect 145 391 146 396
rect 150 391 154 396
rect 158 391 163 396
rect 168 391 169 396
rect 185 391 189 396
rect 194 391 197 396
rect 206 391 207 396
rect 212 391 214 396
rect 218 391 222 396
rect 226 391 227 396
rect 232 391 233 396
rect 237 391 241 396
rect 245 391 250 396
rect 255 391 256 396
rect 11 332 15 337
rect 20 332 23 337
rect 32 332 33 337
rect 38 332 40 337
rect 44 332 48 337
rect 52 332 53 337
rect 58 332 59 337
rect 63 332 67 337
rect 71 332 76 337
rect 81 332 82 337
rect 98 332 102 337
rect 107 332 110 337
rect 119 332 120 337
rect 125 332 127 337
rect 131 332 135 337
rect 139 332 140 337
rect 145 332 146 337
rect 150 332 154 337
rect 158 332 163 337
rect 168 332 169 337
rect 185 332 189 337
rect 194 332 197 337
rect 206 332 207 337
rect 212 332 214 337
rect 218 332 222 337
rect 226 332 227 337
rect 232 332 233 337
rect 237 332 241 337
rect 245 332 250 337
rect 255 332 256 337
rect 11 273 15 278
rect 20 273 23 278
rect 32 273 33 278
rect 38 273 40 278
rect 44 273 48 278
rect 52 273 53 278
rect 58 273 59 278
rect 63 273 67 278
rect 71 273 76 278
rect 81 273 82 278
rect 98 273 102 278
rect 107 273 110 278
rect 119 273 120 278
rect 125 273 127 278
rect 131 273 135 278
rect 139 273 140 278
rect 145 273 146 278
rect 150 273 154 278
rect 158 273 163 278
rect 168 273 169 278
rect 185 273 189 278
rect 194 273 197 278
rect 206 273 207 278
rect 212 273 214 278
rect 218 273 222 278
rect 226 273 227 278
rect 232 273 233 278
rect 237 273 241 278
rect 245 273 250 278
rect 255 273 256 278
rect 11 214 15 219
rect 20 214 23 219
rect 32 214 33 219
rect 38 214 40 219
rect 44 214 48 219
rect 52 214 53 219
rect 58 214 59 219
rect 63 214 67 219
rect 71 214 76 219
rect 81 214 82 219
rect 98 214 102 219
rect 107 214 110 219
rect 119 214 120 219
rect 125 214 127 219
rect 131 214 135 219
rect 139 214 140 219
rect 145 214 146 219
rect 150 214 154 219
rect 158 214 163 219
rect 168 214 169 219
rect 185 214 189 219
rect 194 214 197 219
rect 206 214 207 219
rect 212 214 214 219
rect 218 214 222 219
rect 226 214 227 219
rect 232 214 233 219
rect 237 214 241 219
rect 245 214 250 219
rect 255 214 256 219
rect 11 155 15 160
rect 20 155 23 160
rect 32 155 33 160
rect 38 155 40 160
rect 44 155 48 160
rect 52 155 53 160
rect 58 155 59 160
rect 63 155 67 160
rect 71 155 76 160
rect 81 155 82 160
rect 98 155 102 160
rect 107 155 110 160
rect 119 155 120 160
rect 125 155 127 160
rect 131 155 135 160
rect 139 155 140 160
rect 145 155 146 160
rect 150 155 154 160
rect 158 155 163 160
rect 168 155 169 160
rect 185 155 189 160
rect 194 155 197 160
rect 206 155 207 160
rect 212 155 214 160
rect 218 155 222 160
rect 226 155 227 160
rect 232 155 233 160
rect 237 155 241 160
rect 245 155 250 160
rect 255 155 256 160
rect 11 96 15 101
rect 20 96 23 101
rect 32 96 33 101
rect 38 96 40 101
rect 44 96 48 101
rect 52 96 53 101
rect 58 96 59 101
rect 63 96 67 101
rect 71 96 76 101
rect 81 96 82 101
rect 98 96 102 101
rect 107 96 110 101
rect 119 96 120 101
rect 125 96 127 101
rect 131 96 135 101
rect 139 96 140 101
rect 145 96 146 101
rect 150 96 154 101
rect 158 96 163 101
rect 168 96 169 101
rect 185 96 189 101
rect 194 96 197 101
rect 206 96 207 101
rect 212 96 214 101
rect 218 96 222 101
rect 226 96 227 101
rect 232 96 233 101
rect 237 96 241 101
rect 245 96 250 101
rect 255 96 256 101
rect 11 37 15 42
rect 20 37 23 42
rect 32 37 33 42
rect 38 37 40 42
rect 44 37 48 42
rect 52 37 53 42
rect 58 37 59 42
rect 63 37 67 42
rect 71 37 76 42
rect 81 37 82 42
rect 98 37 102 42
rect 107 37 110 42
rect 119 37 120 42
rect 125 37 127 42
rect 131 37 135 42
rect 139 37 140 42
rect 145 37 146 42
rect 150 37 154 42
rect 158 37 163 42
rect 168 37 169 42
rect 185 37 189 42
rect 194 37 197 42
rect 206 37 207 42
rect 212 37 214 42
rect 218 37 222 42
rect 226 37 227 42
rect 232 37 233 42
rect 237 37 241 42
rect 245 37 250 42
rect 255 37 256 42
<< ndcontact >>
rect 6 433 11 438
rect 23 433 28 438
rect 33 433 38 438
rect 53 433 58 438
rect 76 433 81 438
rect 93 433 98 438
rect 110 433 115 438
rect 120 433 125 438
rect 140 433 145 438
rect 163 433 168 438
rect 180 433 185 438
rect 197 433 202 438
rect 207 433 212 438
rect 227 433 232 438
rect 250 433 255 438
rect 6 374 11 379
rect 23 374 28 379
rect 33 374 38 379
rect 53 374 58 379
rect 76 374 81 379
rect 93 374 98 379
rect 110 374 115 379
rect 120 374 125 379
rect 140 374 145 379
rect 163 374 168 379
rect 180 374 185 379
rect 197 374 202 379
rect 207 374 212 379
rect 227 374 232 379
rect 250 374 255 379
rect 6 315 11 320
rect 23 315 28 320
rect 33 315 38 320
rect 53 315 58 320
rect 76 315 81 320
rect 93 315 98 320
rect 110 315 115 320
rect 120 315 125 320
rect 140 315 145 320
rect 163 315 168 320
rect 180 315 185 320
rect 197 315 202 320
rect 207 315 212 320
rect 227 315 232 320
rect 250 315 255 320
rect 6 256 11 261
rect 23 256 28 261
rect 33 256 38 261
rect 53 256 58 261
rect 76 256 81 261
rect 93 256 98 261
rect 110 256 115 261
rect 120 256 125 261
rect 140 256 145 261
rect 163 256 168 261
rect 180 256 185 261
rect 197 256 202 261
rect 207 256 212 261
rect 227 256 232 261
rect 250 256 255 261
rect 6 197 11 202
rect 23 197 28 202
rect 33 197 38 202
rect 53 197 58 202
rect 76 197 81 202
rect 93 197 98 202
rect 110 197 115 202
rect 120 197 125 202
rect 140 197 145 202
rect 163 197 168 202
rect 180 197 185 202
rect 197 197 202 202
rect 207 197 212 202
rect 227 197 232 202
rect 250 197 255 202
rect 6 138 11 143
rect 23 138 28 143
rect 33 138 38 143
rect 53 138 58 143
rect 76 138 81 143
rect 93 138 98 143
rect 110 138 115 143
rect 120 138 125 143
rect 140 138 145 143
rect 163 138 168 143
rect 180 138 185 143
rect 197 138 202 143
rect 207 138 212 143
rect 227 138 232 143
rect 250 138 255 143
rect 6 79 11 84
rect 23 79 28 84
rect 33 79 38 84
rect 53 79 58 84
rect 76 79 81 84
rect 93 79 98 84
rect 110 79 115 84
rect 120 79 125 84
rect 140 79 145 84
rect 163 79 168 84
rect 180 79 185 84
rect 197 79 202 84
rect 207 79 212 84
rect 227 79 232 84
rect 250 79 255 84
rect 6 20 11 25
rect 23 20 28 25
rect 33 20 38 25
rect 53 20 58 25
rect 76 20 81 25
rect 93 20 98 25
rect 110 20 115 25
rect 120 20 125 25
rect 140 20 145 25
rect 163 20 168 25
rect 180 20 185 25
rect 197 20 202 25
rect 207 20 212 25
rect 227 20 232 25
rect 250 20 255 25
<< pdcontact >>
rect 6 450 11 455
rect 23 450 28 455
rect 33 450 38 455
rect 53 450 58 455
rect 76 450 81 455
rect 93 450 98 455
rect 110 450 115 455
rect 120 450 125 455
rect 140 450 145 455
rect 163 450 168 455
rect 180 450 185 455
rect 197 450 202 455
rect 207 450 212 455
rect 227 450 232 455
rect 250 450 255 455
rect 6 391 11 396
rect 23 391 28 396
rect 33 391 38 396
rect 53 391 58 396
rect 76 391 81 396
rect 93 391 98 396
rect 110 391 115 396
rect 120 391 125 396
rect 140 391 145 396
rect 163 391 168 396
rect 180 391 185 396
rect 197 391 202 396
rect 207 391 212 396
rect 227 391 232 396
rect 250 391 255 396
rect 6 332 11 337
rect 23 332 28 337
rect 33 332 38 337
rect 53 332 58 337
rect 76 332 81 337
rect 93 332 98 337
rect 110 332 115 337
rect 120 332 125 337
rect 140 332 145 337
rect 163 332 168 337
rect 180 332 185 337
rect 197 332 202 337
rect 207 332 212 337
rect 227 332 232 337
rect 250 332 255 337
rect 6 273 11 278
rect 23 273 28 278
rect 33 273 38 278
rect 53 273 58 278
rect 76 273 81 278
rect 93 273 98 278
rect 110 273 115 278
rect 120 273 125 278
rect 140 273 145 278
rect 163 273 168 278
rect 180 273 185 278
rect 197 273 202 278
rect 207 273 212 278
rect 227 273 232 278
rect 250 273 255 278
rect 6 214 11 219
rect 23 214 28 219
rect 33 214 38 219
rect 53 214 58 219
rect 76 214 81 219
rect 93 214 98 219
rect 110 214 115 219
rect 120 214 125 219
rect 140 214 145 219
rect 163 214 168 219
rect 180 214 185 219
rect 197 214 202 219
rect 207 214 212 219
rect 227 214 232 219
rect 250 214 255 219
rect 6 155 11 160
rect 23 155 28 160
rect 33 155 38 160
rect 53 155 58 160
rect 76 155 81 160
rect 93 155 98 160
rect 110 155 115 160
rect 120 155 125 160
rect 140 155 145 160
rect 163 155 168 160
rect 180 155 185 160
rect 197 155 202 160
rect 207 155 212 160
rect 227 155 232 160
rect 250 155 255 160
rect 6 96 11 101
rect 23 96 28 101
rect 33 96 38 101
rect 53 96 58 101
rect 76 96 81 101
rect 93 96 98 101
rect 110 96 115 101
rect 120 96 125 101
rect 140 96 145 101
rect 163 96 168 101
rect 180 96 185 101
rect 197 96 202 101
rect 207 96 212 101
rect 227 96 232 101
rect 250 96 255 101
rect 6 37 11 42
rect 23 37 28 42
rect 33 37 38 42
rect 53 37 58 42
rect 76 37 81 42
rect 93 37 98 42
rect 110 37 115 42
rect 120 37 125 42
rect 140 37 145 42
rect 163 37 168 42
rect 180 37 185 42
rect 197 37 202 42
rect 207 37 212 42
rect 227 37 232 42
rect 250 37 255 42
<< polysilicon >>
rect 15 455 20 459
rect 40 455 44 460
rect 48 455 52 458
rect 59 455 63 458
rect 67 455 71 460
rect 102 455 107 459
rect 127 455 131 460
rect 135 455 139 458
rect 146 455 150 458
rect 154 455 158 460
rect 189 455 194 459
rect 214 455 218 460
rect 222 455 226 458
rect 233 455 237 458
rect 241 455 245 460
rect 15 447 20 450
rect 15 438 20 442
rect 40 438 44 450
rect 48 446 52 450
rect 59 446 63 450
rect 48 438 52 442
rect 59 438 63 442
rect 67 438 71 450
rect 102 447 107 450
rect 102 438 107 442
rect 127 438 131 450
rect 135 446 139 450
rect 146 446 150 450
rect 135 438 139 442
rect 146 438 150 442
rect 154 438 158 450
rect 189 447 194 450
rect 189 438 194 442
rect 214 438 218 450
rect 222 446 226 450
rect 233 446 237 450
rect 222 438 226 442
rect 233 438 237 442
rect 241 438 245 450
rect 15 427 20 433
rect 40 420 44 433
rect 48 430 52 433
rect 59 427 63 433
rect 67 426 71 433
rect 102 427 107 433
rect 127 420 131 433
rect 135 430 139 433
rect 146 427 150 433
rect 154 426 158 433
rect 189 427 194 433
rect 214 420 218 433
rect 222 430 226 433
rect 233 427 237 433
rect 241 426 245 433
rect 15 396 20 400
rect 40 396 44 401
rect 48 396 52 399
rect 59 396 63 399
rect 67 396 71 401
rect 102 396 107 400
rect 127 396 131 401
rect 135 396 139 399
rect 146 396 150 399
rect 154 396 158 401
rect 189 396 194 400
rect 214 396 218 401
rect 222 396 226 399
rect 233 396 237 399
rect 241 396 245 401
rect 15 388 20 391
rect 15 379 20 383
rect 40 379 44 391
rect 48 387 52 391
rect 59 387 63 391
rect 48 379 52 383
rect 59 379 63 383
rect 67 379 71 391
rect 102 388 107 391
rect 102 379 107 383
rect 127 379 131 391
rect 135 387 139 391
rect 146 387 150 391
rect 135 379 139 383
rect 146 379 150 383
rect 154 379 158 391
rect 189 388 194 391
rect 189 379 194 383
rect 214 379 218 391
rect 222 387 226 391
rect 233 387 237 391
rect 222 379 226 383
rect 233 379 237 383
rect 241 379 245 391
rect 15 368 20 374
rect 40 361 44 374
rect 48 371 52 374
rect 59 368 63 374
rect 67 367 71 374
rect 102 368 107 374
rect 127 361 131 374
rect 135 371 139 374
rect 146 368 150 374
rect 154 367 158 374
rect 189 368 194 374
rect 214 361 218 374
rect 222 371 226 374
rect 233 368 237 374
rect 241 367 245 374
rect 15 337 20 341
rect 40 337 44 342
rect 48 337 52 340
rect 59 337 63 340
rect 67 337 71 342
rect 102 337 107 341
rect 127 337 131 342
rect 135 337 139 340
rect 146 337 150 340
rect 154 337 158 342
rect 189 337 194 341
rect 214 337 218 342
rect 222 337 226 340
rect 233 337 237 340
rect 241 337 245 342
rect 15 329 20 332
rect 15 320 20 324
rect 40 320 44 332
rect 48 328 52 332
rect 59 328 63 332
rect 48 320 52 324
rect 59 320 63 324
rect 67 320 71 332
rect 102 329 107 332
rect 102 320 107 324
rect 127 320 131 332
rect 135 328 139 332
rect 146 328 150 332
rect 135 320 139 324
rect 146 320 150 324
rect 154 320 158 332
rect 189 329 194 332
rect 189 320 194 324
rect 214 320 218 332
rect 222 328 226 332
rect 233 328 237 332
rect 222 320 226 324
rect 233 320 237 324
rect 241 320 245 332
rect 15 309 20 315
rect 40 302 44 315
rect 48 312 52 315
rect 59 309 63 315
rect 67 308 71 315
rect 102 309 107 315
rect 127 302 131 315
rect 135 312 139 315
rect 146 309 150 315
rect 154 308 158 315
rect 189 309 194 315
rect 214 302 218 315
rect 222 312 226 315
rect 233 309 237 315
rect 241 308 245 315
rect 15 278 20 282
rect 40 278 44 283
rect 48 278 52 281
rect 59 278 63 281
rect 67 278 71 283
rect 102 278 107 282
rect 127 278 131 283
rect 135 278 139 281
rect 146 278 150 281
rect 154 278 158 283
rect 189 278 194 282
rect 214 278 218 283
rect 222 278 226 281
rect 233 278 237 281
rect 241 278 245 283
rect 15 270 20 273
rect 15 261 20 265
rect 40 261 44 273
rect 48 269 52 273
rect 59 269 63 273
rect 48 261 52 265
rect 59 261 63 265
rect 67 261 71 273
rect 102 270 107 273
rect 102 261 107 265
rect 127 261 131 273
rect 135 269 139 273
rect 146 269 150 273
rect 135 261 139 265
rect 146 261 150 265
rect 154 261 158 273
rect 189 270 194 273
rect 189 261 194 265
rect 214 261 218 273
rect 222 269 226 273
rect 233 269 237 273
rect 222 261 226 265
rect 233 261 237 265
rect 241 261 245 273
rect 15 250 20 256
rect 40 243 44 256
rect 48 253 52 256
rect 59 250 63 256
rect 67 249 71 256
rect 102 250 107 256
rect 127 243 131 256
rect 135 253 139 256
rect 146 250 150 256
rect 154 249 158 256
rect 189 250 194 256
rect 214 243 218 256
rect 222 253 226 256
rect 233 250 237 256
rect 241 249 245 256
rect 15 219 20 223
rect 40 219 44 224
rect 48 219 52 222
rect 59 219 63 222
rect 67 219 71 224
rect 102 219 107 223
rect 127 219 131 224
rect 135 219 139 222
rect 146 219 150 222
rect 154 219 158 224
rect 189 219 194 223
rect 214 219 218 224
rect 222 219 226 222
rect 233 219 237 222
rect 241 219 245 224
rect 15 211 20 214
rect 15 202 20 206
rect 40 202 44 214
rect 48 210 52 214
rect 59 210 63 214
rect 48 202 52 206
rect 59 202 63 206
rect 67 202 71 214
rect 102 211 107 214
rect 102 202 107 206
rect 127 202 131 214
rect 135 210 139 214
rect 146 210 150 214
rect 135 202 139 206
rect 146 202 150 206
rect 154 202 158 214
rect 189 211 194 214
rect 189 202 194 206
rect 214 202 218 214
rect 222 210 226 214
rect 233 210 237 214
rect 222 202 226 206
rect 233 202 237 206
rect 241 202 245 214
rect 15 191 20 197
rect 40 184 44 197
rect 48 194 52 197
rect 59 191 63 197
rect 67 190 71 197
rect 102 191 107 197
rect 127 184 131 197
rect 135 194 139 197
rect 146 191 150 197
rect 154 190 158 197
rect 189 191 194 197
rect 214 184 218 197
rect 222 194 226 197
rect 233 191 237 197
rect 241 190 245 197
rect 15 160 20 164
rect 40 160 44 165
rect 48 160 52 163
rect 59 160 63 163
rect 67 160 71 165
rect 102 160 107 164
rect 127 160 131 165
rect 135 160 139 163
rect 146 160 150 163
rect 154 160 158 165
rect 189 160 194 164
rect 214 160 218 165
rect 222 160 226 163
rect 233 160 237 163
rect 241 160 245 165
rect 15 152 20 155
rect 15 143 20 147
rect 40 143 44 155
rect 48 151 52 155
rect 59 151 63 155
rect 48 143 52 147
rect 59 143 63 147
rect 67 143 71 155
rect 102 152 107 155
rect 102 143 107 147
rect 127 143 131 155
rect 135 151 139 155
rect 146 151 150 155
rect 135 143 139 147
rect 146 143 150 147
rect 154 143 158 155
rect 189 152 194 155
rect 189 143 194 147
rect 214 143 218 155
rect 222 151 226 155
rect 233 151 237 155
rect 222 143 226 147
rect 233 143 237 147
rect 241 143 245 155
rect 15 132 20 138
rect 40 125 44 138
rect 48 135 52 138
rect 59 132 63 138
rect 67 131 71 138
rect 102 132 107 138
rect 127 125 131 138
rect 135 135 139 138
rect 146 132 150 138
rect 154 131 158 138
rect 189 132 194 138
rect 214 125 218 138
rect 222 135 226 138
rect 233 132 237 138
rect 241 131 245 138
rect 15 101 20 105
rect 40 101 44 106
rect 48 101 52 104
rect 59 101 63 104
rect 67 101 71 106
rect 102 101 107 105
rect 127 101 131 106
rect 135 101 139 104
rect 146 101 150 104
rect 154 101 158 106
rect 189 101 194 105
rect 214 101 218 106
rect 222 101 226 104
rect 233 101 237 104
rect 241 101 245 106
rect 15 93 20 96
rect 15 84 20 88
rect 40 84 44 96
rect 48 92 52 96
rect 59 92 63 96
rect 48 84 52 88
rect 59 84 63 88
rect 67 84 71 96
rect 102 93 107 96
rect 102 84 107 88
rect 127 84 131 96
rect 135 92 139 96
rect 146 92 150 96
rect 135 84 139 88
rect 146 84 150 88
rect 154 84 158 96
rect 189 93 194 96
rect 189 84 194 88
rect 214 84 218 96
rect 222 92 226 96
rect 233 92 237 96
rect 222 84 226 88
rect 233 84 237 88
rect 241 84 245 96
rect 15 73 20 79
rect 40 66 44 79
rect 48 76 52 79
rect 59 73 63 79
rect 67 72 71 79
rect 102 73 107 79
rect 127 66 131 79
rect 135 76 139 79
rect 146 73 150 79
rect 154 72 158 79
rect 189 73 194 79
rect 214 66 218 79
rect 222 76 226 79
rect 233 73 237 79
rect 241 72 245 79
rect 15 42 20 46
rect 40 42 44 47
rect 48 42 52 45
rect 59 42 63 45
rect 67 42 71 47
rect 102 42 107 46
rect 127 42 131 47
rect 135 42 139 45
rect 146 42 150 45
rect 154 42 158 47
rect 189 42 194 46
rect 214 42 218 47
rect 222 42 226 45
rect 233 42 237 45
rect 241 42 245 47
rect 15 34 20 37
rect 15 25 20 29
rect 40 25 44 37
rect 48 33 52 37
rect 59 33 63 37
rect 48 25 52 29
rect 59 25 63 29
rect 67 25 71 37
rect 102 34 107 37
rect 102 25 107 29
rect 127 25 131 37
rect 135 33 139 37
rect 146 33 150 37
rect 135 25 139 29
rect 146 25 150 29
rect 154 25 158 37
rect 189 34 194 37
rect 189 25 194 29
rect 214 25 218 37
rect 222 33 226 37
rect 233 33 237 37
rect 222 25 226 29
rect 233 25 237 29
rect 241 25 245 37
rect 15 14 20 20
rect 40 7 44 20
rect 48 17 52 20
rect 59 14 63 20
rect 67 13 71 20
rect 102 14 107 20
rect 127 7 131 20
rect 135 17 139 20
rect 146 14 150 20
rect 154 13 158 20
rect 189 14 194 20
rect 214 7 218 20
rect 222 17 226 20
rect 233 14 237 20
rect 241 13 245 20
<< polycontact >>
rect 48 458 53 463
rect 58 458 63 463
rect 135 458 140 463
rect 145 458 150 463
rect 222 458 227 463
rect 232 458 237 463
rect 15 442 20 447
rect 102 442 107 447
rect 189 442 194 447
rect 48 425 53 430
rect 58 422 63 427
rect 67 421 72 426
rect 135 425 140 430
rect 145 422 150 427
rect 154 421 159 426
rect 222 425 227 430
rect 232 422 237 427
rect 241 421 246 426
rect 39 415 44 420
rect 126 415 131 420
rect 213 415 218 420
rect 48 399 53 404
rect 58 399 63 404
rect 135 399 140 404
rect 145 399 150 404
rect 222 399 227 404
rect 232 399 237 404
rect 15 383 20 388
rect 102 383 107 388
rect 189 383 194 388
rect 48 366 53 371
rect 58 363 63 368
rect 67 362 72 367
rect 135 366 140 371
rect 145 363 150 368
rect 154 362 159 367
rect 222 366 227 371
rect 232 363 237 368
rect 241 362 246 367
rect 39 356 44 361
rect 126 356 131 361
rect 213 356 218 361
rect 48 340 53 345
rect 58 340 63 345
rect 135 340 140 345
rect 145 340 150 345
rect 222 340 227 345
rect 232 340 237 345
rect 15 324 20 329
rect 102 324 107 329
rect 189 324 194 329
rect 48 307 53 312
rect 58 304 63 309
rect 67 303 72 308
rect 135 307 140 312
rect 145 304 150 309
rect 154 303 159 308
rect 222 307 227 312
rect 232 304 237 309
rect 241 303 246 308
rect 39 297 44 302
rect 126 297 131 302
rect 213 297 218 302
rect 48 281 53 286
rect 58 281 63 286
rect 135 281 140 286
rect 145 281 150 286
rect 222 281 227 286
rect 232 281 237 286
rect 15 265 20 270
rect 102 265 107 270
rect 189 265 194 270
rect 48 248 53 253
rect 58 245 63 250
rect 67 244 72 249
rect 135 248 140 253
rect 145 245 150 250
rect 154 244 159 249
rect 222 248 227 253
rect 232 245 237 250
rect 241 244 246 249
rect 39 238 44 243
rect 126 238 131 243
rect 213 238 218 243
rect 48 222 53 227
rect 58 222 63 227
rect 135 222 140 227
rect 145 222 150 227
rect 222 222 227 227
rect 232 222 237 227
rect 15 206 20 211
rect 102 206 107 211
rect 189 206 194 211
rect 48 189 53 194
rect 58 186 63 191
rect 67 185 72 190
rect 135 189 140 194
rect 145 186 150 191
rect 154 185 159 190
rect 222 189 227 194
rect 232 186 237 191
rect 241 185 246 190
rect 39 179 44 184
rect 126 179 131 184
rect 213 179 218 184
rect 48 163 53 168
rect 58 163 63 168
rect 135 163 140 168
rect 145 163 150 168
rect 222 163 227 168
rect 232 163 237 168
rect 15 147 20 152
rect 102 147 107 152
rect 189 147 194 152
rect 48 130 53 135
rect 58 127 63 132
rect 67 126 72 131
rect 135 130 140 135
rect 145 127 150 132
rect 154 126 159 131
rect 222 130 227 135
rect 232 127 237 132
rect 241 126 246 131
rect 39 120 44 125
rect 126 120 131 125
rect 213 120 218 125
rect 48 104 53 109
rect 58 104 63 109
rect 135 104 140 109
rect 145 104 150 109
rect 222 104 227 109
rect 232 104 237 109
rect 15 88 20 93
rect 102 88 107 93
rect 189 88 194 93
rect 48 71 53 76
rect 58 68 63 73
rect 67 67 72 72
rect 135 71 140 76
rect 145 68 150 73
rect 154 67 159 72
rect 222 71 227 76
rect 232 68 237 73
rect 241 67 246 72
rect 39 61 44 66
rect 126 61 131 66
rect 213 61 218 66
rect 48 45 53 50
rect 58 45 63 50
rect 135 45 140 50
rect 145 45 150 50
rect 222 45 227 50
rect 232 45 237 50
rect 15 29 20 34
rect 102 29 107 34
rect 189 29 194 34
rect 48 12 53 17
rect 58 9 63 14
rect 67 8 72 13
rect 135 12 140 17
rect 145 9 150 14
rect 154 8 159 13
rect 222 12 227 17
rect 232 9 237 14
rect 241 8 246 13
rect 39 2 44 7
rect 126 2 131 7
rect 213 2 218 7
<< metal1 >>
rect 50 467 111 470
rect 50 463 53 467
rect 17 460 48 463
rect 5 455 12 456
rect 5 450 6 455
rect 11 450 12 455
rect 5 449 12 450
rect 17 447 20 460
rect 58 463 88 464
rect 107 463 111 467
rect 145 463 175 464
rect 232 463 262 464
rect 63 461 88 463
rect 32 455 39 456
rect 75 455 82 456
rect 5 438 12 439
rect 5 433 6 438
rect 11 433 12 438
rect 5 432 12 433
rect 17 428 20 442
rect 25 438 28 450
rect 32 450 33 455
rect 38 450 39 455
rect 32 449 39 450
rect 54 444 58 450
rect 75 450 76 455
rect 81 450 82 455
rect 75 449 82 450
rect 63 444 70 447
rect 54 441 70 444
rect 25 429 28 433
rect 32 438 39 439
rect 54 438 58 441
rect 63 440 70 441
rect 32 433 33 438
rect 38 433 39 438
rect 75 438 82 439
rect 75 433 76 438
rect 81 433 82 438
rect 32 432 39 433
rect 75 432 82 433
rect 14 421 21 428
rect 25 426 48 429
rect 38 415 39 420
rect 50 417 53 425
rect 57 427 64 428
rect 57 422 58 427
rect 63 422 64 427
rect 57 421 64 422
rect 72 421 73 426
rect 85 417 88 461
rect 104 460 135 463
rect 92 455 99 456
rect 92 450 93 455
rect 98 450 99 455
rect 92 449 99 450
rect 104 447 107 460
rect 150 461 175 463
rect 119 455 126 456
rect 162 455 169 456
rect 92 438 99 439
rect 92 433 93 438
rect 98 433 99 438
rect 92 432 99 433
rect 104 428 107 442
rect 112 438 115 450
rect 119 450 120 455
rect 125 450 126 455
rect 119 449 126 450
rect 141 444 145 450
rect 162 450 163 455
rect 168 450 169 455
rect 162 449 169 450
rect 150 444 157 447
rect 141 441 157 444
rect 112 429 115 433
rect 119 438 126 439
rect 141 438 145 441
rect 150 440 157 441
rect 119 433 120 438
rect 125 433 126 438
rect 162 438 169 439
rect 162 433 163 438
rect 168 433 169 438
rect 119 432 126 433
rect 162 432 169 433
rect 101 421 108 428
rect 112 426 135 429
rect 50 414 88 417
rect 125 415 126 420
rect 137 416 140 425
rect 144 427 151 428
rect 144 422 145 427
rect 150 422 151 427
rect 144 421 151 422
rect 159 421 160 426
rect 172 416 175 461
rect 191 460 222 463
rect 179 455 186 456
rect 179 450 180 455
rect 185 450 186 455
rect 179 449 186 450
rect 191 447 194 460
rect 237 461 262 463
rect 206 455 213 456
rect 249 455 256 456
rect 179 438 186 439
rect 179 433 180 438
rect 185 433 186 438
rect 179 432 186 433
rect 191 428 194 442
rect 199 438 202 450
rect 206 450 207 455
rect 212 450 213 455
rect 206 449 213 450
rect 228 444 232 450
rect 249 450 250 455
rect 255 450 256 455
rect 249 449 256 450
rect 237 444 244 447
rect 228 441 244 444
rect 199 429 202 433
rect 206 438 213 439
rect 228 438 232 441
rect 237 440 244 441
rect 206 433 207 438
rect 212 433 213 438
rect 249 438 256 439
rect 249 433 250 438
rect 255 433 256 438
rect 206 432 213 433
rect 249 432 256 433
rect 188 421 195 428
rect 199 426 222 429
rect 137 413 175 416
rect 212 415 213 420
rect 218 415 219 419
rect 212 412 219 415
rect 224 416 227 425
rect 231 427 238 428
rect 231 422 232 427
rect 237 422 238 427
rect 242 426 250 428
rect 231 421 238 422
rect 246 421 250 426
rect 242 420 250 421
rect 259 416 262 461
rect 224 413 262 416
rect 50 408 111 411
rect 50 404 53 408
rect 17 401 48 404
rect 5 396 12 397
rect 5 391 6 396
rect 11 391 12 396
rect 5 390 12 391
rect 17 388 20 401
rect 58 404 88 405
rect 107 404 111 408
rect 145 404 175 405
rect 232 404 262 405
rect 63 402 88 404
rect 32 396 39 397
rect 75 396 82 397
rect 5 379 12 380
rect 5 374 6 379
rect 11 374 12 379
rect 5 373 12 374
rect 17 369 20 383
rect 25 379 28 391
rect 32 391 33 396
rect 38 391 39 396
rect 32 390 39 391
rect 54 385 58 391
rect 75 391 76 396
rect 81 391 82 396
rect 75 390 82 391
rect 63 385 70 388
rect 54 382 70 385
rect 25 370 28 374
rect 32 379 39 380
rect 54 379 58 382
rect 63 381 70 382
rect 32 374 33 379
rect 38 374 39 379
rect 75 379 82 380
rect 75 374 76 379
rect 81 374 82 379
rect 32 373 39 374
rect 75 373 82 374
rect 14 362 21 369
rect 25 367 48 370
rect 38 356 39 361
rect 50 358 53 366
rect 57 368 64 369
rect 57 363 58 368
rect 63 363 64 368
rect 57 362 64 363
rect 72 362 73 367
rect 85 358 88 402
rect 104 401 135 404
rect 92 396 99 397
rect 92 391 93 396
rect 98 391 99 396
rect 92 390 99 391
rect 104 388 107 401
rect 150 402 175 404
rect 119 396 126 397
rect 162 396 169 397
rect 92 379 99 380
rect 92 374 93 379
rect 98 374 99 379
rect 92 373 99 374
rect 104 369 107 383
rect 112 379 115 391
rect 119 391 120 396
rect 125 391 126 396
rect 119 390 126 391
rect 141 385 145 391
rect 162 391 163 396
rect 168 391 169 396
rect 162 390 169 391
rect 150 385 157 388
rect 141 382 157 385
rect 112 370 115 374
rect 119 379 126 380
rect 141 379 145 382
rect 150 381 157 382
rect 119 374 120 379
rect 125 374 126 379
rect 162 379 169 380
rect 162 374 163 379
rect 168 374 169 379
rect 119 373 126 374
rect 162 373 169 374
rect 101 362 108 369
rect 112 367 135 370
rect 50 355 88 358
rect 125 356 126 361
rect 137 357 140 366
rect 144 368 151 369
rect 144 363 145 368
rect 150 363 151 368
rect 144 362 151 363
rect 159 362 160 367
rect 172 357 175 402
rect 191 401 222 404
rect 179 396 186 397
rect 179 391 180 396
rect 185 391 186 396
rect 179 390 186 391
rect 191 388 194 401
rect 237 402 262 404
rect 206 396 213 397
rect 249 396 256 397
rect 179 379 186 380
rect 179 374 180 379
rect 185 374 186 379
rect 179 373 186 374
rect 191 369 194 383
rect 199 379 202 391
rect 206 391 207 396
rect 212 391 213 396
rect 206 390 213 391
rect 228 385 232 391
rect 249 391 250 396
rect 255 391 256 396
rect 249 390 256 391
rect 237 385 244 388
rect 228 382 244 385
rect 199 370 202 374
rect 206 379 213 380
rect 228 379 232 382
rect 237 381 244 382
rect 206 374 207 379
rect 212 374 213 379
rect 249 379 256 380
rect 249 374 250 379
rect 255 374 256 379
rect 206 373 213 374
rect 249 373 256 374
rect 188 362 195 369
rect 199 367 222 370
rect 137 354 175 357
rect 212 356 213 361
rect 218 356 219 360
rect 212 353 219 356
rect 224 357 227 366
rect 231 368 238 369
rect 231 363 232 368
rect 237 363 238 368
rect 242 367 250 369
rect 231 362 238 363
rect 246 362 250 367
rect 242 361 250 362
rect 259 357 262 402
rect 224 354 262 357
rect 50 349 111 352
rect 50 345 53 349
rect 17 342 48 345
rect 5 337 12 338
rect 5 332 6 337
rect 11 332 12 337
rect 5 331 12 332
rect 17 329 20 342
rect 58 345 88 346
rect 107 345 111 349
rect 145 345 175 346
rect 232 345 262 346
rect 63 343 88 345
rect 32 337 39 338
rect 75 337 82 338
rect 5 320 12 321
rect 5 315 6 320
rect 11 315 12 320
rect 5 314 12 315
rect 17 310 20 324
rect 25 320 28 332
rect 32 332 33 337
rect 38 332 39 337
rect 32 331 39 332
rect 54 326 58 332
rect 75 332 76 337
rect 81 332 82 337
rect 75 331 82 332
rect 63 326 70 329
rect 54 323 70 326
rect 25 311 28 315
rect 32 320 39 321
rect 54 320 58 323
rect 63 322 70 323
rect 32 315 33 320
rect 38 315 39 320
rect 75 320 82 321
rect 75 315 76 320
rect 81 315 82 320
rect 32 314 39 315
rect 75 314 82 315
rect 14 303 21 310
rect 25 308 48 311
rect 38 297 39 302
rect 50 299 53 307
rect 57 309 64 310
rect 57 304 58 309
rect 63 304 64 309
rect 57 303 64 304
rect 72 303 73 308
rect 85 299 88 343
rect 104 342 135 345
rect 92 337 99 338
rect 92 332 93 337
rect 98 332 99 337
rect 92 331 99 332
rect 104 329 107 342
rect 150 343 175 345
rect 119 337 126 338
rect 162 337 169 338
rect 92 320 99 321
rect 92 315 93 320
rect 98 315 99 320
rect 92 314 99 315
rect 104 310 107 324
rect 112 320 115 332
rect 119 332 120 337
rect 125 332 126 337
rect 119 331 126 332
rect 141 326 145 332
rect 162 332 163 337
rect 168 332 169 337
rect 162 331 169 332
rect 150 326 157 329
rect 141 323 157 326
rect 112 311 115 315
rect 119 320 126 321
rect 141 320 145 323
rect 150 322 157 323
rect 119 315 120 320
rect 125 315 126 320
rect 162 320 169 321
rect 162 315 163 320
rect 168 315 169 320
rect 119 314 126 315
rect 162 314 169 315
rect 101 303 108 310
rect 112 308 135 311
rect 50 296 88 299
rect 125 297 126 302
rect 137 298 140 307
rect 144 309 151 310
rect 144 304 145 309
rect 150 304 151 309
rect 144 303 151 304
rect 159 303 160 308
rect 172 298 175 343
rect 191 342 222 345
rect 179 337 186 338
rect 179 332 180 337
rect 185 332 186 337
rect 179 331 186 332
rect 191 329 194 342
rect 237 343 262 345
rect 206 337 213 338
rect 249 337 256 338
rect 179 320 186 321
rect 179 315 180 320
rect 185 315 186 320
rect 179 314 186 315
rect 191 310 194 324
rect 199 320 202 332
rect 206 332 207 337
rect 212 332 213 337
rect 206 331 213 332
rect 228 326 232 332
rect 249 332 250 337
rect 255 332 256 337
rect 249 331 256 332
rect 237 326 244 329
rect 228 323 244 326
rect 199 311 202 315
rect 206 320 213 321
rect 228 320 232 323
rect 237 322 244 323
rect 206 315 207 320
rect 212 315 213 320
rect 249 320 256 321
rect 249 315 250 320
rect 255 315 256 320
rect 206 314 213 315
rect 249 314 256 315
rect 188 303 195 310
rect 199 308 222 311
rect 137 295 175 298
rect 212 297 213 302
rect 218 297 219 301
rect 212 294 219 297
rect 224 298 227 307
rect 231 309 238 310
rect 231 304 232 309
rect 237 304 238 309
rect 242 308 250 310
rect 231 303 238 304
rect 246 303 250 308
rect 242 302 250 303
rect 259 298 262 343
rect 224 295 262 298
rect 50 290 111 293
rect 50 286 53 290
rect 17 283 48 286
rect 5 278 12 279
rect 5 273 6 278
rect 11 273 12 278
rect 5 272 12 273
rect 17 270 20 283
rect 58 286 88 287
rect 107 286 111 290
rect 145 286 175 287
rect 232 286 262 287
rect 63 284 88 286
rect 32 278 39 279
rect 75 278 82 279
rect 5 261 12 262
rect 5 256 6 261
rect 11 256 12 261
rect 5 255 12 256
rect 17 251 20 265
rect 25 261 28 273
rect 32 273 33 278
rect 38 273 39 278
rect 32 272 39 273
rect 54 267 58 273
rect 75 273 76 278
rect 81 273 82 278
rect 75 272 82 273
rect 63 267 70 270
rect 54 264 70 267
rect 25 252 28 256
rect 32 261 39 262
rect 54 261 58 264
rect 63 263 70 264
rect 32 256 33 261
rect 38 256 39 261
rect 75 261 82 262
rect 75 256 76 261
rect 81 256 82 261
rect 32 255 39 256
rect 75 255 82 256
rect 14 244 21 251
rect 25 249 48 252
rect 38 238 39 243
rect 50 240 53 248
rect 57 250 64 251
rect 57 245 58 250
rect 63 245 64 250
rect 57 244 64 245
rect 72 244 73 249
rect 85 240 88 284
rect 104 283 135 286
rect 92 278 99 279
rect 92 273 93 278
rect 98 273 99 278
rect 92 272 99 273
rect 104 270 107 283
rect 150 284 175 286
rect 119 278 126 279
rect 162 278 169 279
rect 92 261 99 262
rect 92 256 93 261
rect 98 256 99 261
rect 92 255 99 256
rect 104 251 107 265
rect 112 261 115 273
rect 119 273 120 278
rect 125 273 126 278
rect 119 272 126 273
rect 141 267 145 273
rect 162 273 163 278
rect 168 273 169 278
rect 162 272 169 273
rect 150 267 157 270
rect 141 264 157 267
rect 112 252 115 256
rect 119 261 126 262
rect 141 261 145 264
rect 150 263 157 264
rect 119 256 120 261
rect 125 256 126 261
rect 162 261 169 262
rect 162 256 163 261
rect 168 256 169 261
rect 119 255 126 256
rect 162 255 169 256
rect 101 244 108 251
rect 112 249 135 252
rect 50 237 88 240
rect 125 238 126 243
rect 137 239 140 248
rect 144 250 151 251
rect 144 245 145 250
rect 150 245 151 250
rect 144 244 151 245
rect 159 244 160 249
rect 172 239 175 284
rect 191 283 222 286
rect 179 278 186 279
rect 179 273 180 278
rect 185 273 186 278
rect 179 272 186 273
rect 191 270 194 283
rect 237 284 262 286
rect 206 278 213 279
rect 249 278 256 279
rect 179 261 186 262
rect 179 256 180 261
rect 185 256 186 261
rect 179 255 186 256
rect 191 251 194 265
rect 199 261 202 273
rect 206 273 207 278
rect 212 273 213 278
rect 206 272 213 273
rect 228 267 232 273
rect 249 273 250 278
rect 255 273 256 278
rect 249 272 256 273
rect 237 267 244 270
rect 228 264 244 267
rect 199 252 202 256
rect 206 261 213 262
rect 228 261 232 264
rect 237 263 244 264
rect 206 256 207 261
rect 212 256 213 261
rect 249 261 256 262
rect 249 256 250 261
rect 255 256 256 261
rect 206 255 213 256
rect 249 255 256 256
rect 188 244 195 251
rect 199 249 222 252
rect 137 236 175 239
rect 212 238 213 243
rect 218 238 219 242
rect 212 235 219 238
rect 224 239 227 248
rect 231 250 238 251
rect 231 245 232 250
rect 237 245 238 250
rect 242 249 250 251
rect 231 244 238 245
rect 246 244 250 249
rect 242 243 250 244
rect 259 239 262 284
rect 224 236 262 239
rect 50 231 111 234
rect 50 227 53 231
rect 17 224 48 227
rect 5 219 12 220
rect 5 214 6 219
rect 11 214 12 219
rect 5 213 12 214
rect 17 211 20 224
rect 58 227 88 228
rect 107 227 111 231
rect 145 227 175 228
rect 232 227 262 228
rect 63 225 88 227
rect 32 219 39 220
rect 75 219 82 220
rect 5 202 12 203
rect 5 197 6 202
rect 11 197 12 202
rect 5 196 12 197
rect 17 192 20 206
rect 25 202 28 214
rect 32 214 33 219
rect 38 214 39 219
rect 32 213 39 214
rect 54 208 58 214
rect 75 214 76 219
rect 81 214 82 219
rect 75 213 82 214
rect 63 208 70 211
rect 54 205 70 208
rect 25 193 28 197
rect 32 202 39 203
rect 54 202 58 205
rect 63 204 70 205
rect 32 197 33 202
rect 38 197 39 202
rect 75 202 82 203
rect 75 197 76 202
rect 81 197 82 202
rect 32 196 39 197
rect 75 196 82 197
rect 14 185 21 192
rect 25 190 48 193
rect 38 179 39 184
rect 50 181 53 189
rect 57 191 64 192
rect 57 186 58 191
rect 63 186 64 191
rect 57 185 64 186
rect 72 185 73 190
rect 85 181 88 225
rect 104 224 135 227
rect 92 219 99 220
rect 92 214 93 219
rect 98 214 99 219
rect 92 213 99 214
rect 104 211 107 224
rect 150 225 175 227
rect 119 219 126 220
rect 162 219 169 220
rect 92 202 99 203
rect 92 197 93 202
rect 98 197 99 202
rect 92 196 99 197
rect 104 192 107 206
rect 112 202 115 214
rect 119 214 120 219
rect 125 214 126 219
rect 119 213 126 214
rect 141 208 145 214
rect 162 214 163 219
rect 168 214 169 219
rect 162 213 169 214
rect 150 208 157 211
rect 141 205 157 208
rect 112 193 115 197
rect 119 202 126 203
rect 141 202 145 205
rect 150 204 157 205
rect 119 197 120 202
rect 125 197 126 202
rect 162 202 169 203
rect 162 197 163 202
rect 168 197 169 202
rect 119 196 126 197
rect 162 196 169 197
rect 101 185 108 192
rect 112 190 135 193
rect 50 178 88 181
rect 125 179 126 184
rect 137 180 140 189
rect 144 191 151 192
rect 144 186 145 191
rect 150 186 151 191
rect 144 185 151 186
rect 159 185 160 190
rect 172 180 175 225
rect 191 224 222 227
rect 179 219 186 220
rect 179 214 180 219
rect 185 214 186 219
rect 179 213 186 214
rect 191 211 194 224
rect 237 225 262 227
rect 206 219 213 220
rect 249 219 256 220
rect 179 202 186 203
rect 179 197 180 202
rect 185 197 186 202
rect 179 196 186 197
rect 191 192 194 206
rect 199 202 202 214
rect 206 214 207 219
rect 212 214 213 219
rect 206 213 213 214
rect 228 208 232 214
rect 249 214 250 219
rect 255 214 256 219
rect 249 213 256 214
rect 237 208 244 211
rect 228 205 244 208
rect 199 193 202 197
rect 206 202 213 203
rect 228 202 232 205
rect 237 204 244 205
rect 206 197 207 202
rect 212 197 213 202
rect 249 202 256 203
rect 249 197 250 202
rect 255 197 256 202
rect 206 196 213 197
rect 249 196 256 197
rect 188 185 195 192
rect 199 190 222 193
rect 137 177 175 180
rect 212 179 213 184
rect 218 179 219 183
rect 212 176 219 179
rect 224 180 227 189
rect 231 191 238 192
rect 231 186 232 191
rect 237 186 238 191
rect 242 190 250 192
rect 231 185 238 186
rect 246 185 250 190
rect 242 184 250 185
rect 259 180 262 225
rect 224 177 262 180
rect 50 172 111 175
rect 50 168 53 172
rect 17 165 48 168
rect 5 160 12 161
rect 5 155 6 160
rect 11 155 12 160
rect 5 154 12 155
rect 17 152 20 165
rect 58 168 88 169
rect 107 168 111 172
rect 145 168 175 169
rect 232 168 262 169
rect 63 166 88 168
rect 32 160 39 161
rect 75 160 82 161
rect 5 143 12 144
rect 5 138 6 143
rect 11 138 12 143
rect 5 137 12 138
rect 17 133 20 147
rect 25 143 28 155
rect 32 155 33 160
rect 38 155 39 160
rect 32 154 39 155
rect 54 149 58 155
rect 75 155 76 160
rect 81 155 82 160
rect 75 154 82 155
rect 63 149 70 152
rect 54 146 70 149
rect 25 134 28 138
rect 32 143 39 144
rect 54 143 58 146
rect 63 145 70 146
rect 32 138 33 143
rect 38 138 39 143
rect 75 143 82 144
rect 75 138 76 143
rect 81 138 82 143
rect 32 137 39 138
rect 75 137 82 138
rect 14 126 21 133
rect 25 131 48 134
rect 38 120 39 125
rect 50 122 53 130
rect 57 132 64 133
rect 57 127 58 132
rect 63 127 64 132
rect 57 126 64 127
rect 72 126 73 131
rect 85 122 88 166
rect 104 165 135 168
rect 92 160 99 161
rect 92 155 93 160
rect 98 155 99 160
rect 92 154 99 155
rect 104 152 107 165
rect 150 166 175 168
rect 119 160 126 161
rect 162 160 169 161
rect 92 143 99 144
rect 92 138 93 143
rect 98 138 99 143
rect 92 137 99 138
rect 104 133 107 147
rect 112 143 115 155
rect 119 155 120 160
rect 125 155 126 160
rect 119 154 126 155
rect 141 149 145 155
rect 162 155 163 160
rect 168 155 169 160
rect 162 154 169 155
rect 150 149 157 152
rect 141 146 157 149
rect 112 134 115 138
rect 119 143 126 144
rect 141 143 145 146
rect 150 145 157 146
rect 119 138 120 143
rect 125 138 126 143
rect 162 143 169 144
rect 162 138 163 143
rect 168 138 169 143
rect 119 137 126 138
rect 162 137 169 138
rect 101 126 108 133
rect 112 131 135 134
rect 50 119 88 122
rect 125 120 126 125
rect 137 121 140 130
rect 144 132 151 133
rect 144 127 145 132
rect 150 127 151 132
rect 144 126 151 127
rect 159 126 160 131
rect 172 121 175 166
rect 191 165 222 168
rect 179 160 186 161
rect 179 155 180 160
rect 185 155 186 160
rect 179 154 186 155
rect 191 152 194 165
rect 237 166 262 168
rect 206 160 213 161
rect 249 160 256 161
rect 179 143 186 144
rect 179 138 180 143
rect 185 138 186 143
rect 179 137 186 138
rect 191 133 194 147
rect 199 143 202 155
rect 206 155 207 160
rect 212 155 213 160
rect 206 154 213 155
rect 228 149 232 155
rect 249 155 250 160
rect 255 155 256 160
rect 249 154 256 155
rect 237 149 244 152
rect 228 146 244 149
rect 199 134 202 138
rect 206 143 213 144
rect 228 143 232 146
rect 237 145 244 146
rect 206 138 207 143
rect 212 138 213 143
rect 249 143 256 144
rect 249 138 250 143
rect 255 138 256 143
rect 206 137 213 138
rect 249 137 256 138
rect 188 126 195 133
rect 199 131 222 134
rect 137 118 175 121
rect 212 120 213 125
rect 218 120 219 124
rect 212 117 219 120
rect 224 121 227 130
rect 231 132 238 133
rect 231 127 232 132
rect 237 127 238 132
rect 242 131 250 133
rect 231 126 238 127
rect 246 126 250 131
rect 242 125 250 126
rect 259 121 262 166
rect 224 118 262 121
rect 50 113 111 116
rect 50 109 53 113
rect 17 106 48 109
rect 5 101 12 102
rect 5 96 6 101
rect 11 96 12 101
rect 5 95 12 96
rect 17 93 20 106
rect 58 109 88 110
rect 107 109 111 113
rect 145 109 175 110
rect 232 109 262 110
rect 63 107 88 109
rect 32 101 39 102
rect 75 101 82 102
rect 5 84 12 85
rect 5 79 6 84
rect 11 79 12 84
rect 5 78 12 79
rect 17 74 20 88
rect 25 84 28 96
rect 32 96 33 101
rect 38 96 39 101
rect 32 95 39 96
rect 54 90 58 96
rect 75 96 76 101
rect 81 96 82 101
rect 75 95 82 96
rect 63 90 70 93
rect 54 87 70 90
rect 25 75 28 79
rect 32 84 39 85
rect 54 84 58 87
rect 63 86 70 87
rect 32 79 33 84
rect 38 79 39 84
rect 75 84 82 85
rect 75 79 76 84
rect 81 79 82 84
rect 32 78 39 79
rect 75 78 82 79
rect 14 67 21 74
rect 25 72 48 75
rect 38 61 39 66
rect 50 63 53 71
rect 57 73 64 74
rect 57 68 58 73
rect 63 68 64 73
rect 57 67 64 68
rect 72 67 73 72
rect 85 63 88 107
rect 104 106 135 109
rect 92 101 99 102
rect 92 96 93 101
rect 98 96 99 101
rect 92 95 99 96
rect 104 93 107 106
rect 150 107 175 109
rect 119 101 126 102
rect 162 101 169 102
rect 92 84 99 85
rect 92 79 93 84
rect 98 79 99 84
rect 92 78 99 79
rect 104 74 107 88
rect 112 84 115 96
rect 119 96 120 101
rect 125 96 126 101
rect 119 95 126 96
rect 141 90 145 96
rect 162 96 163 101
rect 168 96 169 101
rect 162 95 169 96
rect 150 90 157 93
rect 141 87 157 90
rect 112 75 115 79
rect 119 84 126 85
rect 141 84 145 87
rect 150 86 157 87
rect 119 79 120 84
rect 125 79 126 84
rect 162 84 169 85
rect 162 79 163 84
rect 168 79 169 84
rect 119 78 126 79
rect 162 78 169 79
rect 101 67 108 74
rect 112 72 135 75
rect 50 60 88 63
rect 125 61 126 66
rect 137 62 140 71
rect 144 73 151 74
rect 144 68 145 73
rect 150 68 151 73
rect 144 67 151 68
rect 159 67 160 72
rect 172 62 175 107
rect 191 106 222 109
rect 179 101 186 102
rect 179 96 180 101
rect 185 96 186 101
rect 179 95 186 96
rect 191 93 194 106
rect 237 107 262 109
rect 206 101 213 102
rect 249 101 256 102
rect 179 84 186 85
rect 179 79 180 84
rect 185 79 186 84
rect 179 78 186 79
rect 191 74 194 88
rect 199 84 202 96
rect 206 96 207 101
rect 212 96 213 101
rect 206 95 213 96
rect 228 90 232 96
rect 249 96 250 101
rect 255 96 256 101
rect 249 95 256 96
rect 237 90 244 93
rect 228 87 244 90
rect 199 75 202 79
rect 206 84 213 85
rect 228 84 232 87
rect 237 86 244 87
rect 206 79 207 84
rect 212 79 213 84
rect 249 84 256 85
rect 249 79 250 84
rect 255 79 256 84
rect 206 78 213 79
rect 249 78 256 79
rect 188 67 195 74
rect 199 72 222 75
rect 137 59 175 62
rect 212 61 213 66
rect 218 61 219 65
rect 212 58 219 61
rect 224 62 227 71
rect 231 73 238 74
rect 231 68 232 73
rect 237 68 238 73
rect 242 72 250 74
rect 231 67 238 68
rect 246 67 250 72
rect 242 66 250 67
rect 259 62 262 107
rect 224 59 262 62
rect 50 54 111 57
rect 50 50 53 54
rect 17 47 48 50
rect 5 42 12 43
rect 5 37 6 42
rect 11 37 12 42
rect 5 36 12 37
rect 17 34 20 47
rect 58 50 88 51
rect 107 50 111 54
rect 145 50 175 51
rect 232 50 262 51
rect 63 48 88 50
rect 32 42 39 43
rect 75 42 82 43
rect 5 25 12 26
rect 5 20 6 25
rect 11 20 12 25
rect 5 19 12 20
rect 17 15 20 29
rect 25 25 28 37
rect 32 37 33 42
rect 38 37 39 42
rect 32 36 39 37
rect 54 31 58 37
rect 75 37 76 42
rect 81 37 82 42
rect 75 36 82 37
rect 63 31 70 34
rect 54 28 70 31
rect 25 16 28 20
rect 32 25 39 26
rect 54 25 58 28
rect 63 27 70 28
rect 32 20 33 25
rect 38 20 39 25
rect 75 25 82 26
rect 75 20 76 25
rect 81 20 82 25
rect 32 19 39 20
rect 75 19 82 20
rect 14 8 21 15
rect 25 13 48 16
rect 38 2 39 7
rect 50 4 53 12
rect 57 14 64 15
rect 57 9 58 14
rect 63 9 64 14
rect 57 8 64 9
rect 72 8 73 13
rect 85 4 88 48
rect 104 47 135 50
rect 92 42 99 43
rect 92 37 93 42
rect 98 37 99 42
rect 92 36 99 37
rect 104 34 107 47
rect 150 48 175 50
rect 119 42 126 43
rect 162 42 169 43
rect 92 25 99 26
rect 92 20 93 25
rect 98 20 99 25
rect 92 19 99 20
rect 104 15 107 29
rect 112 25 115 37
rect 119 37 120 42
rect 125 37 126 42
rect 119 36 126 37
rect 141 31 145 37
rect 162 37 163 42
rect 168 37 169 42
rect 162 36 169 37
rect 150 31 157 34
rect 141 28 157 31
rect 112 16 115 20
rect 119 25 126 26
rect 141 25 145 28
rect 150 27 157 28
rect 119 20 120 25
rect 125 20 126 25
rect 162 25 169 26
rect 162 20 163 25
rect 168 20 169 25
rect 119 19 126 20
rect 162 19 169 20
rect 101 8 108 15
rect 112 13 135 16
rect 50 1 88 4
rect 125 2 126 7
rect 137 3 140 12
rect 144 14 151 15
rect 144 9 145 14
rect 150 9 151 14
rect 144 8 151 9
rect 159 8 160 13
rect 172 3 175 48
rect 191 47 222 50
rect 179 42 186 43
rect 179 37 180 42
rect 185 37 186 42
rect 179 36 186 37
rect 191 34 194 47
rect 237 48 262 50
rect 206 42 213 43
rect 249 42 256 43
rect 179 25 186 26
rect 179 20 180 25
rect 185 20 186 25
rect 179 19 186 20
rect 191 15 194 29
rect 199 25 202 37
rect 206 37 207 42
rect 212 37 213 42
rect 206 36 213 37
rect 228 31 232 37
rect 249 37 250 42
rect 255 37 256 42
rect 249 36 256 37
rect 237 31 244 34
rect 228 28 244 31
rect 199 16 202 20
rect 206 25 213 26
rect 228 25 232 28
rect 237 27 244 28
rect 206 20 207 25
rect 212 20 213 25
rect 249 25 256 26
rect 249 20 250 25
rect 255 20 256 25
rect 206 19 213 20
rect 249 19 256 20
rect 188 8 195 15
rect 199 13 222 16
rect 137 0 175 3
rect 212 2 213 7
rect 218 2 219 6
rect 212 -1 219 2
rect 224 3 227 12
rect 231 14 238 15
rect 231 9 232 14
rect 237 9 238 14
rect 242 13 250 15
rect 231 8 238 9
rect 246 8 250 13
rect 242 7 250 8
rect 259 3 262 48
rect 224 0 262 3
<< metal2 >>
rect -2 455 1 470
rect 5 455 12 456
rect 32 455 39 456
rect 75 455 82 456
rect 92 455 99 456
rect 119 455 126 456
rect 162 455 169 456
rect 179 455 186 456
rect 206 455 213 456
rect 249 455 256 456
rect -2 451 256 455
rect -2 450 58 451
rect -2 396 1 450
rect 5 449 12 450
rect 32 449 39 450
rect 75 449 82 451
rect 92 450 145 451
rect 162 450 232 451
rect 92 449 99 450
rect 119 449 126 450
rect 162 449 169 450
rect 179 449 186 450
rect 206 449 213 450
rect 249 449 256 451
rect 63 440 70 447
rect 150 440 157 447
rect 237 440 244 447
rect 5 438 12 439
rect 32 438 39 439
rect 5 436 58 438
rect 75 437 82 439
rect 92 438 99 439
rect 119 438 126 439
rect 92 437 145 438
rect 75 436 145 437
rect 162 437 169 439
rect 179 438 186 439
rect 206 438 213 439
rect 249 438 256 439
rect 260 438 263 470
rect 179 437 232 438
rect 162 436 232 437
rect 249 436 263 438
rect 5 433 263 436
rect 5 432 12 433
rect 32 432 39 433
rect 75 432 82 433
rect 92 432 99 433
rect 119 432 126 433
rect 162 432 169 433
rect 179 432 186 433
rect 206 432 213 433
rect 249 432 256 433
rect 14 427 21 428
rect 57 427 64 428
rect 14 423 64 427
rect 14 421 21 423
rect 57 421 64 423
rect 101 427 108 428
rect 144 427 151 428
rect 101 423 151 427
rect 101 421 108 423
rect 144 421 151 423
rect 188 427 195 428
rect 231 427 238 428
rect 188 423 238 427
rect 188 421 195 423
rect 231 421 238 423
rect 242 420 250 428
rect 212 412 219 419
rect 5 396 12 397
rect 32 396 39 397
rect 75 396 82 397
rect 92 396 99 397
rect 119 396 126 397
rect 162 396 169 397
rect 179 396 186 397
rect 206 396 213 397
rect 249 396 256 397
rect -2 392 256 396
rect -2 391 58 392
rect -2 337 1 391
rect 5 390 12 391
rect 32 390 39 391
rect 75 390 82 392
rect 92 391 145 392
rect 162 391 232 392
rect 92 390 99 391
rect 119 390 126 391
rect 162 390 169 391
rect 179 390 186 391
rect 206 390 213 391
rect 249 390 256 392
rect 63 381 70 388
rect 150 381 157 388
rect 237 381 244 388
rect 5 379 12 380
rect 32 379 39 380
rect 5 377 58 379
rect 75 378 82 380
rect 92 379 99 380
rect 119 379 126 380
rect 92 378 145 379
rect 75 377 145 378
rect 162 378 169 380
rect 179 379 186 380
rect 206 379 213 380
rect 249 379 256 380
rect 260 379 263 433
rect 179 378 232 379
rect 162 377 232 378
rect 249 377 263 379
rect 5 374 263 377
rect 5 373 12 374
rect 32 373 39 374
rect 75 373 82 374
rect 92 373 99 374
rect 119 373 126 374
rect 162 373 169 374
rect 179 373 186 374
rect 206 373 213 374
rect 249 373 256 374
rect 14 368 21 369
rect 57 368 64 369
rect 14 364 64 368
rect 14 362 21 364
rect 57 362 64 364
rect 101 368 108 369
rect 144 368 151 369
rect 101 364 151 368
rect 101 362 108 364
rect 144 362 151 364
rect 188 368 195 369
rect 231 368 238 369
rect 188 364 238 368
rect 188 362 195 364
rect 231 362 238 364
rect 242 361 250 369
rect 212 353 219 360
rect 5 337 12 338
rect 32 337 39 338
rect 75 337 82 338
rect 92 337 99 338
rect 119 337 126 338
rect 162 337 169 338
rect 179 337 186 338
rect 206 337 213 338
rect 249 337 256 338
rect -2 333 256 337
rect -2 332 58 333
rect -2 278 1 332
rect 5 331 12 332
rect 32 331 39 332
rect 75 331 82 333
rect 92 332 145 333
rect 162 332 232 333
rect 92 331 99 332
rect 119 331 126 332
rect 162 331 169 332
rect 179 331 186 332
rect 206 331 213 332
rect 249 331 256 333
rect 63 322 70 329
rect 150 322 157 329
rect 237 322 244 329
rect 5 320 12 321
rect 32 320 39 321
rect 5 318 58 320
rect 75 319 82 321
rect 92 320 99 321
rect 119 320 126 321
rect 92 319 145 320
rect 75 318 145 319
rect 162 319 169 321
rect 179 320 186 321
rect 206 320 213 321
rect 249 320 256 321
rect 260 320 263 374
rect 179 319 232 320
rect 162 318 232 319
rect 249 318 263 320
rect 5 315 263 318
rect 5 314 12 315
rect 32 314 39 315
rect 75 314 82 315
rect 92 314 99 315
rect 119 314 126 315
rect 162 314 169 315
rect 179 314 186 315
rect 206 314 213 315
rect 249 314 256 315
rect 14 309 21 310
rect 57 309 64 310
rect 14 305 64 309
rect 14 303 21 305
rect 57 303 64 305
rect 101 309 108 310
rect 144 309 151 310
rect 101 305 151 309
rect 101 303 108 305
rect 144 303 151 305
rect 188 309 195 310
rect 231 309 238 310
rect 188 305 238 309
rect 188 303 195 305
rect 231 303 238 305
rect 242 302 250 310
rect 212 294 219 301
rect 5 278 12 279
rect 32 278 39 279
rect 75 278 82 279
rect 92 278 99 279
rect 119 278 126 279
rect 162 278 169 279
rect 179 278 186 279
rect 206 278 213 279
rect 249 278 256 279
rect -2 274 256 278
rect -2 273 58 274
rect -2 219 1 273
rect 5 272 12 273
rect 32 272 39 273
rect 75 272 82 274
rect 92 273 145 274
rect 162 273 232 274
rect 92 272 99 273
rect 119 272 126 273
rect 162 272 169 273
rect 179 272 186 273
rect 206 272 213 273
rect 249 272 256 274
rect 63 263 70 270
rect 150 263 157 270
rect 237 263 244 270
rect 5 261 12 262
rect 32 261 39 262
rect 5 259 58 261
rect 75 260 82 262
rect 92 261 99 262
rect 119 261 126 262
rect 92 260 145 261
rect 75 259 145 260
rect 162 260 169 262
rect 179 261 186 262
rect 206 261 213 262
rect 249 261 256 262
rect 260 261 263 315
rect 179 260 232 261
rect 162 259 232 260
rect 249 259 263 261
rect 5 256 263 259
rect 5 255 12 256
rect 32 255 39 256
rect 75 255 82 256
rect 92 255 99 256
rect 119 255 126 256
rect 162 255 169 256
rect 179 255 186 256
rect 206 255 213 256
rect 249 255 256 256
rect 14 250 21 251
rect 57 250 64 251
rect 14 246 64 250
rect 14 244 21 246
rect 57 244 64 246
rect 101 250 108 251
rect 144 250 151 251
rect 101 246 151 250
rect 101 244 108 246
rect 144 244 151 246
rect 188 250 195 251
rect 231 250 238 251
rect 188 246 238 250
rect 188 244 195 246
rect 231 244 238 246
rect 242 243 250 251
rect 212 235 219 242
rect 5 219 12 220
rect 32 219 39 220
rect 75 219 82 220
rect 92 219 99 220
rect 119 219 126 220
rect 162 219 169 220
rect 179 219 186 220
rect 206 219 213 220
rect 249 219 256 220
rect -2 215 256 219
rect -2 214 58 215
rect -2 160 1 214
rect 5 213 12 214
rect 32 213 39 214
rect 75 213 82 215
rect 92 214 145 215
rect 162 214 232 215
rect 92 213 99 214
rect 119 213 126 214
rect 162 213 169 214
rect 179 213 186 214
rect 206 213 213 214
rect 249 213 256 215
rect 63 204 70 211
rect 150 204 157 211
rect 237 204 244 211
rect 5 202 12 203
rect 32 202 39 203
rect 5 200 58 202
rect 75 201 82 203
rect 92 202 99 203
rect 119 202 126 203
rect 92 201 145 202
rect 75 200 145 201
rect 162 201 169 203
rect 179 202 186 203
rect 206 202 213 203
rect 249 202 256 203
rect 260 202 263 256
rect 179 201 232 202
rect 162 200 232 201
rect 249 200 263 202
rect 5 197 263 200
rect 5 196 12 197
rect 32 196 39 197
rect 75 196 82 197
rect 92 196 99 197
rect 119 196 126 197
rect 162 196 169 197
rect 179 196 186 197
rect 206 196 213 197
rect 249 196 256 197
rect 14 191 21 192
rect 57 191 64 192
rect 14 187 64 191
rect 14 185 21 187
rect 57 185 64 187
rect 101 191 108 192
rect 144 191 151 192
rect 101 187 151 191
rect 101 185 108 187
rect 144 185 151 187
rect 188 191 195 192
rect 231 191 238 192
rect 188 187 238 191
rect 188 185 195 187
rect 231 185 238 187
rect 242 184 250 192
rect 212 176 219 183
rect 5 160 12 161
rect 32 160 39 161
rect 75 160 82 161
rect 92 160 99 161
rect 119 160 126 161
rect 162 160 169 161
rect 179 160 186 161
rect 206 160 213 161
rect 249 160 256 161
rect -2 156 256 160
rect -2 155 58 156
rect -2 101 1 155
rect 5 154 12 155
rect 32 154 39 155
rect 75 154 82 156
rect 92 155 145 156
rect 162 155 232 156
rect 92 154 99 155
rect 119 154 126 155
rect 162 154 169 155
rect 179 154 186 155
rect 206 154 213 155
rect 249 154 256 156
rect 63 145 70 152
rect 150 145 157 152
rect 237 145 244 152
rect 5 143 12 144
rect 32 143 39 144
rect 5 141 58 143
rect 75 142 82 144
rect 92 143 99 144
rect 119 143 126 144
rect 92 142 145 143
rect 75 141 145 142
rect 162 142 169 144
rect 179 143 186 144
rect 206 143 213 144
rect 249 143 256 144
rect 260 143 263 197
rect 179 142 232 143
rect 162 141 232 142
rect 249 141 263 143
rect 5 138 263 141
rect 5 137 12 138
rect 32 137 39 138
rect 75 137 82 138
rect 92 137 99 138
rect 119 137 126 138
rect 162 137 169 138
rect 179 137 186 138
rect 206 137 213 138
rect 249 137 256 138
rect 14 132 21 133
rect 57 132 64 133
rect 14 128 64 132
rect 14 126 21 128
rect 57 126 64 128
rect 101 132 108 133
rect 144 132 151 133
rect 101 128 151 132
rect 101 126 108 128
rect 144 126 151 128
rect 188 132 195 133
rect 231 132 238 133
rect 188 128 238 132
rect 188 126 195 128
rect 231 126 238 128
rect 242 125 250 133
rect 212 117 219 124
rect 5 101 12 102
rect 32 101 39 102
rect 75 101 82 102
rect 92 101 99 102
rect 119 101 126 102
rect 162 101 169 102
rect 179 101 186 102
rect 206 101 213 102
rect 249 101 256 102
rect -2 97 256 101
rect -2 96 58 97
rect -2 42 1 96
rect 5 95 12 96
rect 32 95 39 96
rect 75 95 82 97
rect 92 96 145 97
rect 162 96 232 97
rect 92 95 99 96
rect 119 95 126 96
rect 162 95 169 96
rect 179 95 186 96
rect 206 95 213 96
rect 249 95 256 97
rect 63 86 70 93
rect 150 86 157 93
rect 237 86 244 93
rect 5 84 12 85
rect 32 84 39 85
rect 5 82 58 84
rect 75 83 82 85
rect 92 84 99 85
rect 119 84 126 85
rect 92 83 145 84
rect 75 82 145 83
rect 162 83 169 85
rect 179 84 186 85
rect 206 84 213 85
rect 249 84 256 85
rect 260 84 263 138
rect 179 83 232 84
rect 162 82 232 83
rect 249 82 263 84
rect 5 79 263 82
rect 5 78 12 79
rect 32 78 39 79
rect 75 78 82 79
rect 92 78 99 79
rect 119 78 126 79
rect 162 78 169 79
rect 179 78 186 79
rect 206 78 213 79
rect 249 78 256 79
rect 14 73 21 74
rect 57 73 64 74
rect 14 69 64 73
rect 14 67 21 69
rect 57 67 64 69
rect 101 73 108 74
rect 144 73 151 74
rect 101 69 151 73
rect 101 67 108 69
rect 144 67 151 69
rect 188 73 195 74
rect 231 73 238 74
rect 188 69 238 73
rect 188 67 195 69
rect 231 67 238 69
rect 242 66 250 74
rect 212 58 219 65
rect 5 42 12 43
rect 32 42 39 43
rect 75 42 82 43
rect 92 42 99 43
rect 119 42 126 43
rect 162 42 169 43
rect 179 42 186 43
rect 206 42 213 43
rect 249 42 256 43
rect -2 38 256 42
rect -2 37 58 38
rect -2 -2 1 37
rect 5 36 12 37
rect 32 36 39 37
rect 75 36 82 38
rect 92 37 145 38
rect 162 37 232 38
rect 92 36 99 37
rect 119 36 126 37
rect 162 36 169 37
rect 179 36 186 37
rect 206 36 213 37
rect 249 36 256 38
rect 63 27 70 34
rect 150 27 157 34
rect 237 27 244 34
rect 5 25 12 26
rect 32 25 39 26
rect 5 23 58 25
rect 75 24 82 26
rect 92 25 99 26
rect 119 25 126 26
rect 92 24 145 25
rect 75 23 145 24
rect 162 24 169 26
rect 179 25 186 26
rect 206 25 213 26
rect 249 25 256 26
rect 260 25 263 79
rect 179 24 232 25
rect 162 23 232 24
rect 249 23 263 25
rect 5 20 263 23
rect 5 19 12 20
rect 32 19 39 20
rect 75 19 82 20
rect 92 19 99 20
rect 119 19 126 20
rect 162 19 169 20
rect 179 19 186 20
rect 206 19 213 20
rect 249 19 256 20
rect 14 14 21 15
rect 57 14 64 15
rect 14 10 64 14
rect 14 8 21 10
rect 57 8 64 10
rect 101 14 108 15
rect 144 14 151 15
rect 101 10 151 14
rect 101 8 108 10
rect 144 8 151 10
rect 188 14 195 15
rect 231 14 238 15
rect 188 10 238 14
rect 188 8 195 10
rect 231 8 238 10
rect 242 7 250 15
rect 212 -1 219 6
rect 260 -2 263 20
<< gv1 >>
rect 6 450 11 455
rect 33 450 38 455
rect 76 450 81 455
rect 93 450 98 455
rect 120 450 125 455
rect 163 450 168 455
rect 180 450 185 455
rect 207 450 212 455
rect 250 450 255 455
rect 64 441 69 446
rect 151 441 156 446
rect 238 441 243 446
rect 6 433 11 438
rect 33 433 38 438
rect 76 433 81 438
rect 93 433 98 438
rect 120 433 125 438
rect 163 433 168 438
rect 180 433 185 438
rect 207 433 212 438
rect 250 433 255 438
rect 15 422 20 427
rect 58 422 63 427
rect 102 422 107 427
rect 145 422 150 427
rect 189 422 194 427
rect 232 422 237 427
rect 243 421 249 427
rect 213 413 218 418
rect 6 391 11 396
rect 33 391 38 396
rect 76 391 81 396
rect 93 391 98 396
rect 120 391 125 396
rect 163 391 168 396
rect 180 391 185 396
rect 207 391 212 396
rect 250 391 255 396
rect 64 382 69 387
rect 151 382 156 387
rect 238 382 243 387
rect 6 374 11 379
rect 33 374 38 379
rect 76 374 81 379
rect 93 374 98 379
rect 120 374 125 379
rect 163 374 168 379
rect 180 374 185 379
rect 207 374 212 379
rect 250 374 255 379
rect 15 363 20 368
rect 58 363 63 368
rect 102 363 107 368
rect 145 363 150 368
rect 189 363 194 368
rect 232 363 237 368
rect 243 362 249 368
rect 213 354 218 359
rect 6 332 11 337
rect 33 332 38 337
rect 76 332 81 337
rect 93 332 98 337
rect 120 332 125 337
rect 163 332 168 337
rect 180 332 185 337
rect 207 332 212 337
rect 250 332 255 337
rect 64 323 69 328
rect 151 323 156 328
rect 238 323 243 328
rect 6 315 11 320
rect 33 315 38 320
rect 76 315 81 320
rect 93 315 98 320
rect 120 315 125 320
rect 163 315 168 320
rect 180 315 185 320
rect 207 315 212 320
rect 250 315 255 320
rect 15 304 20 309
rect 58 304 63 309
rect 102 304 107 309
rect 145 304 150 309
rect 189 304 194 309
rect 232 304 237 309
rect 243 303 249 309
rect 213 295 218 300
rect 6 273 11 278
rect 33 273 38 278
rect 76 273 81 278
rect 93 273 98 278
rect 120 273 125 278
rect 163 273 168 278
rect 180 273 185 278
rect 207 273 212 278
rect 250 273 255 278
rect 64 264 69 269
rect 151 264 156 269
rect 238 264 243 269
rect 6 256 11 261
rect 33 256 38 261
rect 76 256 81 261
rect 93 256 98 261
rect 120 256 125 261
rect 163 256 168 261
rect 180 256 185 261
rect 207 256 212 261
rect 250 256 255 261
rect 15 245 20 250
rect 58 245 63 250
rect 102 245 107 250
rect 145 245 150 250
rect 189 245 194 250
rect 232 245 237 250
rect 243 244 249 250
rect 213 236 218 241
rect 6 214 11 219
rect 33 214 38 219
rect 76 214 81 219
rect 93 214 98 219
rect 120 214 125 219
rect 163 214 168 219
rect 180 214 185 219
rect 207 214 212 219
rect 250 214 255 219
rect 64 205 69 210
rect 151 205 156 210
rect 238 205 243 210
rect 6 197 11 202
rect 33 197 38 202
rect 76 197 81 202
rect 93 197 98 202
rect 120 197 125 202
rect 163 197 168 202
rect 180 197 185 202
rect 207 197 212 202
rect 250 197 255 202
rect 15 186 20 191
rect 58 186 63 191
rect 102 186 107 191
rect 145 186 150 191
rect 189 186 194 191
rect 232 186 237 191
rect 243 185 249 191
rect 213 177 218 182
rect 6 155 11 160
rect 33 155 38 160
rect 76 155 81 160
rect 93 155 98 160
rect 120 155 125 160
rect 163 155 168 160
rect 180 155 185 160
rect 207 155 212 160
rect 250 155 255 160
rect 64 146 69 151
rect 151 146 156 151
rect 238 146 243 151
rect 6 138 11 143
rect 33 138 38 143
rect 76 138 81 143
rect 93 138 98 143
rect 120 138 125 143
rect 163 138 168 143
rect 180 138 185 143
rect 207 138 212 143
rect 250 138 255 143
rect 15 127 20 132
rect 58 127 63 132
rect 102 127 107 132
rect 145 127 150 132
rect 189 127 194 132
rect 232 127 237 132
rect 243 126 249 132
rect 213 118 218 123
rect 6 96 11 101
rect 33 96 38 101
rect 76 96 81 101
rect 93 96 98 101
rect 120 96 125 101
rect 163 96 168 101
rect 180 96 185 101
rect 207 96 212 101
rect 250 96 255 101
rect 64 87 69 92
rect 151 87 156 92
rect 238 87 243 92
rect 6 79 11 84
rect 33 79 38 84
rect 76 79 81 84
rect 93 79 98 84
rect 120 79 125 84
rect 163 79 168 84
rect 180 79 185 84
rect 207 79 212 84
rect 250 79 255 84
rect 15 68 20 73
rect 58 68 63 73
rect 102 68 107 73
rect 145 68 150 73
rect 189 68 194 73
rect 232 68 237 73
rect 243 67 249 73
rect 213 59 218 64
rect 6 37 11 42
rect 33 37 38 42
rect 76 37 81 42
rect 93 37 98 42
rect 120 37 125 42
rect 163 37 168 42
rect 180 37 185 42
rect 207 37 212 42
rect 250 37 255 42
rect 64 28 69 33
rect 151 28 156 33
rect 238 28 243 33
rect 6 20 11 25
rect 33 20 38 25
rect 76 20 81 25
rect 93 20 98 25
rect 120 20 125 25
rect 163 20 168 25
rect 180 20 185 25
rect 207 20 212 25
rect 250 20 255 25
rect 15 9 20 14
rect 58 9 63 14
rect 102 9 107 14
rect 145 9 150 14
rect 189 9 194 14
rect 232 9 237 14
rect 243 8 249 14
rect 213 0 218 5
<< metal3 >>
rect 15 428 18 470
rect 63 440 70 447
rect 150 445 157 447
rect 150 441 226 445
rect 150 440 157 441
rect 14 421 21 428
rect 15 369 18 421
rect 64 417 69 440
rect 188 421 195 428
rect 223 425 226 441
rect 242 425 250 428
rect 223 422 250 425
rect 242 420 250 422
rect 212 417 219 419
rect 64 414 219 417
rect 137 413 219 414
rect 212 412 219 413
rect 63 381 70 388
rect 150 386 157 388
rect 150 382 226 386
rect 150 381 157 382
rect 14 362 21 369
rect 15 310 18 362
rect 64 358 69 381
rect 188 362 195 369
rect 223 366 226 382
rect 242 366 250 369
rect 223 363 250 366
rect 242 361 250 363
rect 212 358 219 360
rect 64 355 219 358
rect 137 354 219 355
rect 212 353 219 354
rect 63 322 70 329
rect 150 327 157 329
rect 150 323 226 327
rect 150 322 157 323
rect 14 303 21 310
rect 15 251 18 303
rect 64 299 69 322
rect 188 303 195 310
rect 223 307 226 323
rect 242 307 250 310
rect 223 304 250 307
rect 242 302 250 304
rect 212 299 219 301
rect 64 296 219 299
rect 137 295 219 296
rect 212 294 219 295
rect 63 263 70 270
rect 150 268 157 270
rect 150 264 226 268
rect 150 263 157 264
rect 14 244 21 251
rect 15 192 18 244
rect 64 240 69 263
rect 188 244 195 251
rect 223 248 226 264
rect 242 248 250 251
rect 223 245 250 248
rect 242 243 250 245
rect 212 240 219 242
rect 64 237 219 240
rect 137 236 219 237
rect 212 235 219 236
rect 63 204 70 211
rect 150 209 157 211
rect 150 205 226 209
rect 150 204 157 205
rect 14 185 21 192
rect 15 133 18 185
rect 64 181 69 204
rect 188 185 195 192
rect 223 189 226 205
rect 242 189 250 192
rect 223 186 250 189
rect 242 184 250 186
rect 212 181 219 183
rect 64 178 219 181
rect 137 177 219 178
rect 212 176 219 177
rect 63 145 70 152
rect 150 150 157 152
rect 150 146 226 150
rect 150 145 157 146
rect 14 126 21 133
rect 15 74 18 126
rect 64 122 69 145
rect 188 126 195 133
rect 223 130 226 146
rect 242 130 250 133
rect 223 127 250 130
rect 242 125 250 127
rect 212 122 219 124
rect 64 119 219 122
rect 137 118 219 119
rect 212 117 219 118
rect 63 86 70 93
rect 150 91 157 93
rect 150 87 226 91
rect 150 86 157 87
rect 14 67 21 74
rect 15 15 18 67
rect 64 63 69 86
rect 188 67 195 74
rect 223 71 226 87
rect 242 71 250 74
rect 223 68 250 71
rect 242 66 250 68
rect 212 63 219 65
rect 64 60 219 63
rect 137 59 219 60
rect 212 58 219 59
rect 63 27 70 34
rect 150 32 157 34
rect 150 28 226 32
rect 150 27 157 28
rect 14 8 21 15
rect 15 -2 18 8
rect 64 4 69 27
rect 188 8 195 15
rect 223 12 226 28
rect 242 12 250 15
rect 223 9 250 12
rect 242 7 250 9
rect 212 4 219 6
rect 64 1 219 4
rect 137 0 219 1
rect 212 -1 219 0
<< gv2 >>
rect 64 441 69 446
rect 151 441 156 446
rect 15 422 20 427
rect 189 422 194 427
rect 243 421 249 427
rect 213 413 218 418
rect 64 382 69 387
rect 151 382 156 387
rect 15 363 20 368
rect 189 363 194 368
rect 243 362 249 368
rect 213 354 218 359
rect 64 323 69 328
rect 151 323 156 328
rect 15 304 20 309
rect 189 304 194 309
rect 243 303 249 309
rect 213 295 218 300
rect 64 264 69 269
rect 151 264 156 269
rect 15 245 20 250
rect 189 245 194 250
rect 243 244 249 250
rect 213 236 218 241
rect 64 205 69 210
rect 151 205 156 210
rect 15 186 20 191
rect 189 186 194 191
rect 243 185 249 191
rect 213 177 218 182
rect 64 146 69 151
rect 151 146 156 151
rect 15 127 20 132
rect 189 127 194 132
rect 243 126 249 132
rect 213 118 218 123
rect 64 87 69 92
rect 151 87 156 92
rect 15 68 20 73
rect 189 68 194 73
rect 243 67 249 73
rect 213 59 218 64
rect 64 28 69 33
rect 151 28 156 33
rect 15 9 20 14
rect 189 9 194 14
rect 243 8 249 14
rect 213 0 218 5
<< metal4 >>
rect 190 428 193 470
rect 188 421 195 428
rect 190 369 193 421
rect 188 362 195 369
rect 190 310 193 362
rect 188 303 195 310
rect 190 251 193 303
rect 188 244 195 251
rect 190 192 193 244
rect 188 185 195 192
rect 190 133 193 185
rect 188 126 195 133
rect 190 74 193 126
rect 188 67 195 74
rect 190 15 193 67
rect 188 8 195 15
rect 190 -2 193 8
<< gv3 >>
rect 189 422 194 427
rect 189 363 194 368
rect 189 304 194 309
rect 189 245 194 250
rect 189 186 194 191
rect 189 127 194 132
rect 189 68 194 73
rect 189 9 194 14
<< labels >>
rlabel metal2 -1 38 0 40 3 Vdd!
rlabel metal2 261 23 262 25 7 GND!
rlabel metal3 16 2 17 4 1 b
rlabel metal4 191 5 192 7 1 a
rlabel polycontact 41 4 42 5 1 g0_0
rlabel polycontact 41 63 42 64 1 g0_1
rlabel polycontact 41 122 42 123 1 g0_2
rlabel polycontact 41 181 42 182 1 g0_3
rlabel polycontact 41 240 42 241 1 g0_4
rlabel polycontact 41 299 42 300 1 g0_5
rlabel polycontact 41 358 42 359 1 g0_6
rlabel polycontact 40 416 43 420 1 g0_7
rlabel polycontact 70 424 71 425 1 g1_7
rlabel polycontact 71 364 72 365 1 g1_6
rlabel polycontact 71 305 72 306 1 g1_5
rlabel polycontact 71 245 72 246 1 g1_4
rlabel polycontact 70 187 71 188 1 g1_3
rlabel polycontact 71 128 72 129 1 g1_2
rlabel polycontact 71 68 72 69 1 g1_1
rlabel polycontact 71 9 72 10 1 g1_0
rlabel polycontact 128 5 129 6 1 g2_0
rlabel polycontact 128 65 129 66 1 g2_1
rlabel polycontact 128 123 129 124 1 g2_2
rlabel polycontact 128 183 129 184 1 g2_3
rlabel polycontact 129 241 130 242 1 g2_4
rlabel polycontact 129 301 130 302 1 g2_5
rlabel polycontact 129 359 130 360 1 g2_6
rlabel polycontact 128 418 129 419 1 g2_7
rlabel polycontact 156 10 157 11 1 g3_0
rlabel polycontact 156 69 157 70 1 g3_1
rlabel polycontact 157 128 158 129 1 g3_2
rlabel polycontact 156 186 157 187 1 g3_3
rlabel polycontact 157 246 158 247 1 g3_4
rlabel polycontact 156 305 157 306 1 g3_5
rlabel polycontact 156 364 157 365 1 g3_6
rlabel polycontact 156 422 157 423 1 g3_7
rlabel gv1 239 89 240 90 1 out01
rlabel gv1 239 30 240 31 1 out00
rlabel gv1 240 265 241 266 1 out04
rlabel gv1 240 325 241 326 1 out05
rlabel gv1 238 384 239 385 1 out06
rlabel gv1 238 443 239 444 1 out07
rlabel gv1 238 147 239 148 1 out02
rlabel gv1 238 206 241 208 1 out03
<< end >>
